PK   *�4Wku��"  Gb    cirkitFile.json�ݎ�H��_����d&|7����L7���AP��\�T���h_f�i3X��$�'Yq��L_�������!�b�϶�/�m��l���~{����^H�����_��?uW�w��v�i�v���^��g�����|�w��&�i�~�
}�Y�X����̺eWg}S��2�*�ֵn�����+�Y��bf�*�673X\[��
��f��kCTx�n�k�Ͷ��&9��w��n�����l�̻SwGw��ٸ;�yw*s�X\[��
�m��u�y�ns���Z��bQ�,Ty�y�WY=/��|�bQ5�խ��y����p���ҙ��1� N;����#�3�Y"R��=f�Ha?��%"����.)�N-v�Haw{��S�4S�_;�U"^�گ�����f�H�j�{gn�N�D������#/�s��v6K8�P2S�W Ϲ�3��������f�Hawq�D,��.n��b�Z��3Ba?#�%"�N���Pد������f�Hawq�D����Y"R�}�,)�>l�p����Y"Rد�����f�Ha�N�D� ��{��{�Y"Rؽ�,)��i��v�4KD
�w�%\��i��v�4KD
�w�%"��;����f�Ha�N�D��{�Y"Rؽ�,)��i��v�4K���{�Y"Rؽ�,)��9�0?4`�a�O0�`���m�d�o09;���v�����,M)�}���B�c#�c�J'X:�����A�K�l�<6vP:���S�����gp*�Y*`�>�3�"�%6g��g���h=GA�L�{fT��{��Y(�`�\[ccWcc�,�kl�l�t���gC����z�'`>}2?h� `>��3����+,����i`p����O�|�38~�
�'`>}?p���0�>;���^�|�ӧ���WX>�������+,���t�8~���'`>]#���?�|�������,���t]
8~�oV�_���\����'`��R�w��7~O��˗���� ��/9�|��	�O�\��._�|���^����,���t�8~���'`>]b��|��	�O��-�/X>��J���HY!��뱻'Gv�.p�S��,���t�(8~�g��������K._�|�������,���t�18~���'`>]%��|��	�O�w��._�|�ӕ�����,���tM=6~\�`�̧� �����0��1 �\`�̧���X>�i�p���[�\����\`�̧�:���X>�i�p����O�|�#?p���0�vw�\`�̧}i�����'`>������	�O{���?�|��.F����,�����8~���'`>��z�<z�<����#��,����[8~���'`>�3�����	�O;����?�|���n������'`>�J�����	�O����?�|r�ﱛ�J�Ԯ.��_��y��n�P��t}��Go��8�����m'?��:q�a�Չ���N~��t������6�8��#�Դ���1�Fo��:ޘy���M:�d���R�Upu楮��\��Y��\V������᧣�4�t𓆟�}��A\V�}���Z���"��5�<��������Ջ��E��y��ë*k|��W}����ՙߞ4���OG>i���'?��I�O�|���~�4���&?�I�O�mZ�X�Θwg�6m�1���m��3��ҳ�L��Zچ�	~��3�O~&�)Í�?sԧ?sԧ?sԧ?s�'��5�yw�Oo̼sG}�xc��M�7Z-(��������5��n{���������6�bs���^��(ƣt�on�ov�|!A	9=�`�@BNOa"��ӳ"�$��D�!	�k!��w�ى��T!��?~�mD%��B�H��E�$���V�&X�>
�*�C^���r�h�8���6̷f�(%7\V��`�-0�F)�����o�����pmb�y��L��KoHI;�.,a>��|���`L0�a>�Rzǁ.ys���0G)i�2S����a>�R�VZ0&���0G)i�'X9��BP�f����(%��c��x�G)i_��������	�	����QJڧ��q�q�����1�|��|��}`L�{⸛�0�0G)�w��=��QJ�6��q�q���!F1��t].�	����(%]?
c��x��8JI�9`>`>�R��x0&������t��	��%��QJ��	����㧔�?�u����}i����*GX��0V�.���~d�9��aED�p�\��V�����}\W�PXc�E��asL�Ba=j:o6��D`�
V���\x�b��VDۃ�U���`
�kۆ�U�qe�
�յ��D���2X�ª�s
N�E��>�̉-���ph�mNl9��V8���9'���B+Z}f�[NF��>�ω-�
��
�V�0pb˨n�C+Z]���-���
�Vהpb˩�(�¡յ1��r�2
�phu��N]F���U�ĖS�Qh�C�k�8�%}#F�J�S�场,��eZ���8�89�.;B��EƖS�场�B+Z]�ȉ-�.��
�V�Vrb˩�(�¡�5���r�2
�phu�+'����B+Z]��y0�S�Qh�C�k�9��<�H��c�� p겂S�Qh�C�k�9�%=�Hz\�S����
N]F�����ĖS�Qh�C�=8���eZ��j�Nl9u�V8���[N]F�����ĖS�Qh�C�=8(�����B+Z�%-��2
�ph�'
'����B+Z��-�.��
�V{�pbKZIFZJƩ�<�.󜺌B+Z�ĉ-�.��
�V{qb˩�(�¡�N��r�2
�ph�'����B+Z�E�m��eZ��jo0Nl9u�V8���[N]F���j�ĖS�Qh�C�=�8���eZ��j�<NlI]>Hm>8uY��e�S�Qh�C��9���eZ��jOFNl9u�V8��[�[N]F���ȤĶ��eZ��j�ONl9u�V8�ڳ�[N]F��4��wL�$H��2k�U�y��l�!u�J�WN���{�'���M;Q�D7ى*'�xOT9�y{�ʉ^�UNt���r��D��'����<5�@ɋ��S/}�*���S�V�*s1�e���R�Upu楮��\��Y��\V���	.��rq��T.NS���Y꼸"���o���uV;��||�~�.�%I�b\\�XHYT��w��RUY�k��ݼ��/ŭ.�$�`X.�Q���9JR�x %�\<��T.�	�T.�	�T.�	�T.�	Ҳ����|&H�����3A����r�(\�<���T�)���~Z5��	.��ry�RT.OS���YJQ�<I)*�9��2)*�]&E�ˤ�\v���%/&{\&I��	.�$��`Rx��s�̐�� Se�$^��`����e���à��6�ݮ����u��F����m������r��C�@Bn8[@�@Bn8�@�@Bn8�A�@Bn8#B�@Bn8�B�@Bn8SC�@Bn8�C�@Bn���������"q���m�o̸QJ����n��7J�=\b�`�-0G)��U��f�(%�p	�a��x�q���4�1ᮿq�0�a>�R�ޓ0&���0G)i�C��s�������	��9��QJ��V��|���8JI{���pwRp�R`>^�|��=�`L0/`>�RҞB0&��0G)i��=��QJ�3��q�q����1���n��|��|���`L0�0G)��}��=��QJ�V������QJ�6��� �q�����1���}�	�� �q���Y�1�|<�|��k�`L0/a>�R�5Y0&���0?�4}}�h�Z�a@U(�Bau�h�ZW�PX];Z��Vƕ�*V׎z��U�qe�
�5�]���ڨ@"�`
k���u�B�PX�5
%���)�0X����Q��*0�V���v�7�
�+�U(���LA���`
�>�)8�V8��l3'����Tvq�.�^©�(�¡�g�9��T_Z���3��r*0
�ph��Nl9U�V8����[N%F�����ĖS�Qh�C�kJ8��TdZ����Nl9U�V8��Ƈ���.��
�V�*qb˩�(�¡�5W�ؒ�#}%Ʃ�rN]�s�2
�phu'����B+Z]�ǉ-�.��
�V�$rb˩�(�¡յ���r�2
�phu�('����B+Z]�ʉ-�.��
�V��rL��eZ����cNl9u�V8����[N]F����Ė��"�qEN]Vp겂S�Qh�C�k�9���eZ��j�Nl9u�V8��+�[N]F���|�ĖS�Qh�C��+8���eZ��jJl=�.��
�V{�pb˩�(�¡՞(��r�2
�ph��'����B+Z�QÉ-i%i)�.��s�2
�ph�g'����B+Z�}ĉ-�.��
�V{8qb˩�(�¡�^T��r�2
�ph��%��S�Qh�C���8���eZ��j�3Nl9u�V8�ګ�[N]F�����ĖS�Qh�C���8�%u� ����e�S�N]F���2�ĖS�Qh�C�=9���eZ��joINl9u�V8��#�ےS�Qh�C��>9���eZ��j�RNl9u�V�h��� ��ˬ�Wy�}��[�,ԡ*]_9��S�a��r�7�D��d'����=Q�D��*'zeOT9��z�ʉ~�UNt���r���Ԭ%/&{O��u�&O�Zu�����+K�V�ՙ����s)�fQ.sY-V�'�L���yJR�8MI*g��� .�羉�^�Y��*�E�k�y��$��qq�b!eQe~�-�JUe��}Vv�ϗ���̒��a�8GI*�(I�⁔�r�8JR�x&HR�x&HR�x&HR�x&H�:P�b��� M����i2�38,�ŢpY���jSu��h�>�i�,|W'�L���yJQ�<M)*�g)E��$��`��ˤ�\v���.��r�e������Mp�$L�&�L�&��§�q?U��{o��p��ۮ]ln6�v��m��_�~]o����M������l��v�����_:�-/�S�g����(���&:�i�qѢM�pѝM���}�"�j&2��$��O�9��6i�}�\�P*�;@cTp�j��4��n2^�o=T
�M�a������ ~w��Yq7�\n<�{;}͉��xct��cw�&�~T�������m�v�K�,�n�Ǯ�_F����ן�?�t6p|q��$��x�s|��x���� ;L쯌�h�e����
���oa��w D��_>F�� D�[ ��A�� ν`wH|�@g>��H���q|�3�5�=�D��,�@����:�՗>���K_E��/|��+6,�)s#RoE�1���M{��v����oV�����6��z9{�����A��v�,ᆧ��f	7<�e�0K��)1#�Y�O�)�nxJ���'6�`�*�P���CU��2K��<#�Y���LP�AQt��u$Ya�'X� �خ��y�r �X ~l�pO]Z9 ,f���{x���0^8�]�=<yj�0k�kL�r ?�~j���c8 ~��Ԯ1ܕ�~M���AҊ�W��p7��q�:�xє�֮�/�p �6��]C_N�Yn[�8�*#�|���5�}Q ����Y�����p��v}��`��^��� �^=�^��> �O=�O��� �^-�f-�O=�O��k��S�S���pp ���Ԯ����v�� �i ��]C�38 ~ ~j�о� �����5��,���v�S
� �i	�S����p ����Xü���W���܍�2�����������?�P������׸��Χ8=H:b�����['pz��a���p�F��0�/�O�|��2#�2>�;z��q�G�8=H8G/���=������׸��wD�� ��0�kG���A��0�kG�z��A��0�>���F�+`BA�Ü�bk A
�PDE�]��	M�Ѣc��U���&���1D�+`BA������0��	��kt�W��&4�>4��!�:
�PxG�]��	M��c��R���&ԅ����:L(hB]$��!�N
�Px�c�>��
�N��uJ��S���&��8��Ʀ�	)�l� tZ��0��	���`b�.[���&��W���0��	u�:��L(hB]���!�l
�PW졟A�-`BA�JA�~gojn*h`9l� ��)�U�PЄ��C��a�G��UL����@�-`BA��Zt�e�PЄ�2Ct�&4��jF�]��	M�+��1D�-`BA�jrt�e�PЄ�C�.[���&�U����m
�P;�c��S���&��	���0��	��:��U,�e,�:ţ���S���&Ԏ���0��	�[:��:L(hB�t��!�N
�P���c��S���&�3�t�&4�v�A�]��	M��}�1D�)`BAjW"t�u
�PЄ�Q	Ct�&4�v�B�����]�t��u
�PЄڅCt�&4�vC�]��	M����1D�)`BAj�6pKt�&4�v�C�]��	M���1D�)`B�D���Ε�]]fM��3����2d�U���Iݏ��8q������n�Ǐ��N?�:q��K����Ǐ��N?�&:q�����1'�5�o{�*`����զ
��BY.�b��l\�y��l>�"k�2��b%�YHf�Ɵ����gf��� .�羉�Z�Y�o.�E�k�y�9��I��쿫)�*��n�WU���ge7��|�Kq�s�?i�������3�O� H&��Ɵq��g\8i�Nƅ��ǜ��<��i�<��i�0����&!������ e��HnR�[��RƟs����\ e�9H�sZ3�$	Xs�$	X�P������Uc=oѫ�z��w�������Qg�lw�6��X>���\�^���;#�S��C� �N+��-[�iC�F�6�-E7�Vt�8����.@ǿ.L�r|��e�;�2;�_����n/: ���8��S{��tf�����?���]�y��ex^��L��4�6���I�k���3��Q~������=��f�_��1]0љ^�b���J�� ��G�jc���.��WƄ�)f���t TF9\Am��B����m��t��F=ylƳ?��o��Ǟ8|$�����Ǐ�����0����Q9����Q=����Q1����Q�W��M�$���զ�Y��tΒBZm��u{��?���_�4�����?�]��?�q�y�ow�^/���#d�[on�Y��k'1�Õ��k׸����EEM��1UU7y��z]��y�|�tJ�x׻�.#�Eٮ�]<�I�4��m���=����-���M�q'^f�ϯ#�k���������ɏ�䨼99*�O�*O�
�G�	��
ޟگ���Q�u��������pzTq|��a�������_�7�w3+�r���HR�޾��?4��w���V]�{���O�f�t7������L�/�t�o��ſݽ�����G�ًUws�������w��M��g������>��.=�`x��ޯ���~�o�!<���w������PLM�ʪ��eu��dY~q���l��
}Wf}��YW�L�<kd�̋�*�"�IELʁ����0��{w=�u�4S��Fʲ.�'��4��'c�g%�_����?����^'��>��qJ��Ib���̧N���c�˿t�?k�箚x��Ƀ��q߈�N���鷇<y������q�G����w:wCv�?r�����������zF8���#���o����V�|��.���n��r2��U�������$��*�#�|rV�U���]Wd.�Y]�z)V�W�z���O*�S�����x/����(�|���e��ޯw�|���1��󢼎��O+�U��u(�{�^��d^��Xe���Y��<[�ˏ�6����N�˓��/	y2dC�\L�2z��]]|�A��Y�����`;�u��k�O�M���Q_���?�G�郦:�A.�q�i�?��~_���Q��F�g�j_d��s����2\�}i�*\U�����\���i2x_ǉ�5�^���"Z��Ϻx�[6�>,Fɐrw,1��c�JU��}J�˛U�jG�jF�sl������8�nV���z��������¹I��ijE�Z8Pk�oV���V�;�J'R?ُl^��8H9��w��sd3�����/�tkջ��t���'�Y���x�e�Y��}�ٯ���:��ٛ~��ݲ��k/p����p��{��B�x�/��\v���w�������x�.�޿�.s�پ��x5���*�$ܫ�իx�붻׷�/��,����v	Q��An����E���~�ş'�����^��*��m>h�۬ow?v�7���W�^��>������+�;�鋗���*�sƵE����-�6��o�9w>o��ëه�I�Y��w��Ȭpm8���X�������O͑��㼆��}��r�����fǳD���zp���,ٿg�˒�%G�'gI�4���5'����جt0˙��4��$�y+0}��NL��iܿ�z�;�9��:�j��y�����o>y��\����FNy��f��ן7����$h|,r8	����e�8t4�K�2�Tr��~�t"F���Is=G|G�K���r����4	�YRϒ��ܜ��t��I��c��\�By�X?��L�,���R�͋�U��_$�,9?1M��)��w*|���ݵ����?u�~��ntyï������nﻛo7o���o����ه�PK   Є4WUo�H̒ �� /   images/448c166d-0905-4b6c-8bbe-acf1d9153e5c.png�XUP@����w� A�Cpw� �����=���Kpww]��u�p�zU=3��05U��Ʉ+ȉ##�!   dI	%  R  �����)��@�� ����N�%P�B�B @],"��_o'��  b�g Y8 �g�������E����Ç�ê��E���+���#ÚR��V^pAQ�p|���Ot8{��ʉ���cǣ�MW}�CD���'+��l.ǣ�Iw��쵲�oD4e/���U0�" "�c.,�asrp�`cb.��P��[d����Y���X���-$�\\T�����&���)�4�ߨ�Y�iI�t���s�<��c�)�� L��VVYI��Z����qf��V���j�GGj�
���ɽ�|5_j-*���*���j�ﭻ�%�8ؗL5Ĝ��~�*'��u��ׄD!��Y��p.'%'��~�{U�S嘞������YU�/p§�����r���0�UW3*��� ��;���]Ϋ�DAz�����������c��7;��|��M&,}#���.i�e�o�?�@ |糤��q	ؠ��'X�ꄣ�̔�{S
������?�׼���oB~���,0(x�(���!|H,`%,I��w�����f���)�}u�9���P )��.nnVK_��L���'o�f,,o�*�QH��y��O؏�~qa�1jXJ�PZ*�C�P�^\�ܭG�ӡwR��_��{�����z�᫬�D�2�sR��X8��M�K:����1TTl�g�1�61)�1��3yֹ���	��SS������s�L�OU320�M��XX���r�@�}�r6$mm#'W0��_�(䞐uK�hO�L��lEDF�'0�����!z��Nf��C��+=��{���%�����I֣&� �$��<R�Ӕ[I0F1��虢���u��K,����w�H��`[��R��������zhfJ�lK<<K�TF]*p�2�BZiy���XM\\M��፬9�f�\J\z�|I��P����������,i�}c��ٹaq�����|���!�Y:qmvS ����;�;SqDU�\���6�J�s�Cf?9��S�H��N�A���xP�W�<��r�� %�� �)/[Uތ�]S?��j���m���VJ�S:DC�L�"pM���`te&��YA18 <�q #�]�@71>�Ŀ`����~���	k��ݎ�)��mL�HB�b/�#�J;ј�W?zr?9�����I�mP;IcS�x�+9vf�|�K�q��YC�sr'����RGNm72�n3	�@}�^��l��=�~�/.�2Eh�9���ԣ�җ�w�J����Ƭ���BU�GP�|�U�g2W�srݦ���4ǽ��7<=�o
��s���	_=$A�Ť�� ��pk��SvGr�J+�TX���֖�V��&���i��;��d�1R����<�Q�bE�x,��t*#�nP�Əq3+�q:ƫ4������ �H�5����(���X��ʄ���Z��xrVL���S�3��F�v�ǓYB�ֲF'aQ��c�$�1ᝡ��˄	���*'㱞@�/$��^���Wih�Y�}�d�IN��_�BJ��(����O�?�0kG�^��	���]�K��7�dQAH��R�ս���c � r��].	�������߯�c{'���(��'`�$�3o���%�فq�]~� �"
)]�b3��Ql�i�ɩq�+Y��hr?F�Q��EUv5��&1�j�Z!�9ʸ��T�u�[���1�o�qV�8�NW�;�-���C]��ofl��k�9n:m��pq���[}� g9�*f[?s���&w��%�TM����I���k��G;��r*�	գ�:t�7�mA1����3%%��~մcj�8����pէ��m�zq���VTR���=,+n9�W�GRT�v��`0�!#-m�N��I�S���f
[Y:���7��q��-�k�3��U�h,�h�RPE��X�Lg�4�js�Y
��W���(�KZ.��`5��)ai���S��9}�ro��&�&��؏��+��{���-�
����Kj��Je#�5��K����rU!gƼ�-�1���X�G~<�0o��͟�BH�&h|2"�z4ޑk �i��	�R�@P�8a��������.����&le_)27Q���Qݦ���ǭ<Ƞ���>Y�7��ea����<{����&c�R�P�ciH�M�qJi4c���<�&_\Rq9���d�Y|��������7���p�Ne	�x^6	xo��Dp(�&�91�1�dE�Cn��*�x�"��X���{�����y�x�J��ǵ�6�vl��(�������5*r.��d/�r$�竧"6cR��M�m����� rs��c���̬���@0��AEy�c��,V2?I���xb��D
S(�eb����	]�[�R�T�\��[�h��G3����A4��S������
�':�Kt����V��C��6�^�܏��B����ɢ���b����.���W����Aj?@?��Q[����x�r����蔧|�F��wa�̺������;4jjr-���k�Ze�vG���D���M
����D9�E���K�/�*כN�l*��n�TY��9���Fʈ	䱰�yX=,AɗU��KI�Q�����&�Iz�J����T�Z�	�ٻ�{9�-����f�ە�s�{p|~#ȡ�S���8K�S�B��~�Ѧ��f��l��*��26ظ��ID�����T�UF�:1�����w���D�� ��gh�L/s�_;·{˫��r��%��O���_�5Z��-T�c����"&i1��g��[t�T���	�MK=���*J�Ct`q@@����P�2�^��|�dj�l�!�� ��H��P���FT��4�@���X$�"�г��<	�~��n
p�^�
��e��R�ʟ�Z��ʩ�*��rǥ�vY��K��t]\r�|���L):cb�nKْNV�[l�W锝�ܓ����U�XT^Y0{$]V�	��p+���"`3K�ٙ�����X���5�m����5!�`�]B65]K87z�$��`���C�V��LZ"��t���<�=�h�T��e;4>f��HJ�]^�/�"(��(�.�<l��kmud dDP�r�XQ�C�ޞ�f����8�k�~��wK�6�Y�4G�5���{;��L��݆dj��a����ꋩ��?WGr�x���R
<���6+~��-����a�
��
�&��|kl�߹�����j#ƥ*�K��ʲ�ݳL�C���Nzd�(^7��V�^b??�[��3��N�t7��g�~r"���9���7n <��g����!�������=)ϧ�t���`��Od8(��p4�QU�2�*���EL�}��O�51$��7�D�;j~��X��`��6�������c#ZZXhgt:][D0�b�j\�!E��J;�����>k7SU߿��s�`��Ꜽ�&㛨��p�Dic�O0+tBAȣ�P�$���%�ϓfA���i�'巵�T^kHʁX6��&��.Kp>�|
M�i��̭�ǟ0~~��g�Mj�P�a��z��ʯ�����C}/u]-C���+��͈gL�D=D�F|�~&�8�g��$0�1�Z_��� ��0����u>���r!�te�6/H����,jiHOLH`[=�����2~C�vm������tw璋W%]��g%�ǉ�uF�L����%�|�>�V�0v�*��L��scȦ��c��dC��#Q�f�Q�HF�*~�������	שGW(���4��7��ٓ�mYA\��rôE���¤z��KU`��O�v& VH)�'+�R�<��=a��w;N���lQ�'��P�?
�6�Y+x��ԟ��H��(��J�u_n}|#h�����LH��� ��g��-c�wAuLΏ�B���u�ʸ�]
T�X:	 :?H�_MK�,�C��E����a<]h�+����:��$w^��+{M��3�6J<# �/v,�A7zC%ċ��>��&�V쮯��q�f��W*����8�����<ҹ^�;'�	��(��W"ǐ����zL>q.|�(�����{ai�7K����_\��=:%�������$*Sڭ�bc΃cl�!|�A�2FX.��$�CxCn}�kUb��N𠟿�O�� �u�O�9K,o��7�L�݄��f�4�u���Һ�i�8=�W�Z3;�Z���<����ZY��ƃ����M�� �~yJ�+'%�5��/R���Wv�������N�C� 5��a�#��}b��D���r����?�bo�QIGaT�xGV��M��s���탄Z?�����H#�C�E�;v���-KS�h����C��Ԏ�Y:�jɤ�̡����ʞ�\Y�o�k���W��"��C�i\�.�a0hD�Q��h\"೼��>8�kr��6>,
�k�sr��v�'G��'q��fP~���5��R�����z،�!��e���$�0ݘ�F���
!bz��,��\�=�@��E��i*��db�k7XA��>�k�۬}�l�O��*k*�1��d� 6 �����/�da�J�Y4�H��c)7F�!�ռ�D0�A�^�b��>s�/p|@g���h��xFI��X�y�s���@vAH�i�E���S��NLC/=��Ɂ�0?��j�����m�5����)Qvz��� ьN�	��0�'��d��p�э�`k�~��6w����v*��c�� ��[1 ����e�ۤu�u?��ݖ��=Ű�֡ӧ�AX'3� ��K�r/gB`���0�⫸J�*l�;d�)R�_|��n�I�``�]9U�Y��X�ُ�;:T%�YӚ^���xH�$��2�����<_�9�.��r�bL���p��IqJ�!��͐ዋI=92&��Y���V��J����	�]PP�L~��N�eZ�l�?�w���
��j�JUD�TU�c���#k�߰��rm�)�v&Ms}*������`<����n�B��O:2

���9�h��zk�)����7)")� ٨��R�l�ƹsKJi��J���%GXS$`�|������W�nU�r���d�h�.(�M�����7O�AW?p���7u�/7��f6}8�0�LE���.!��K��U�8�uM��6^,ç����r��%���P����z3�
O�y;#�zy�i��~^i���`c%���0�����<[��-Y�n�q���fˑ.8��)^D4Y.(t��n���{X^K��ˮ�]������0D¤�O8"8��?n		wor�� ���V��v���}x�FT�b�n�!^���	�9�Cy�0_��=3i7O�PNå��������Q� �4+<us���|��.�v�ؿ�=>.�;'�w�'�'�pW�K�=��tC �]�c�Gs��"��6�)���]��fc����l��g�M�x��'>o�74�XC��1u"���?�ڷ^g��lz�9Y�܇��~;�kEqq��n���.:6�{k��V�"/�81��&�+�9�)I���6�����)|-'g����Q
(��)�YA�[�8aƽV��,a�g<Q���	��|��������\�Fv
��hF���c垓�#������w���^/��	�8�e���'D�v}��I��V���y��3WbW{I�z��������i�` <�L8�B*�`;�n���@�tc�<Xy՜,�ڿ]��V�Q	`G""��db���Oi�N �x�B@o{���bRv������S�v���Yl��%(���� ��n���*�Ai����V8g�nW�=}UӃ�+:1=3�.N�����d�ʮ����ѡ�����h����@�:�V��p��$�M� Ǡ֡�H�S�c�m�Z-0+P����f���؛��'w� �8��"�x���ia<D�̹��w[>�Z����q�q��=�Wϧ+���R�/�ʸe�'����JJ�m
q�I�<Ģ�x�p�Y��\���l(m�����*�>V�1�nT���*/i��Cć揄������h7���3�ܥ5U5��e�&"kw.}�N~�x�	Z*��_d��y�_/���':TTՏ�	؜�IC	8l�Of��T%/��-�	0w}~�@�}|���6�k�����b��7��}�(&�0��:�j��%�*}��	�B�>����C7d�_��,�����	9*ݒ�`�ra&��F�zɯ!f��	�Zx����()�_��L �Ć���yϓ��F8CpnA��V4�me�U�t�a�nYv�VUem�y'J�=��`R�Ԕj$��10R�T�r������ �0נ�0H�Y��D�=�b��_�	Rh�+��}L�,��
Z{j�މ��a5Fzf6IN0}��N����ƽMMC��'��Wf$H�֠O"��UO���{p�syW���Y��~�ç{�X���ʂ�*����䶪�;�8��JV�\ �M"�z�M �9P\�!]Ѥ���ӟ(i�<�a��#s���`��ҙ5l�0���m?d'���1�w�G�J0�cZ
�����=s<�L�V-R�a�)���Do�"^��*�f�'W���O"���~�`��zx��}!L�C�'��f��#0�Y*��'Q�vS �+=7?�rja��������3e�$s��ؽ!�sh��~��V������	��o���\]2�ԣd��/#w+�P]HiPV��80��,Sѡ�AX�Ap�͟�r&e���«&w��w�N���� ����R�<�Fz��#	���s�����4�[��.'����nC-���8�xP�T�1������}Vz�������x�ԛ����[}/�+9=DVF`Ru�i�}O�{��ָ�B�|����[����,�?a� ,/I�6^%�%�s�@p�����B=/at��+#� �+���H����I�_��**.护�����o,M����-�-�T�V��]i�$��2͢u��|�mo�?�9�X��g����H�b'`�����S�!�3�`Ukʅ��t��Y� ݪJ��$%�]=n[�t�b=T-i*=��F�\A���{�d,���W<��\|u*�lqze�-Q�DOy9��KPe!w�W������K!W�#�l��G%3��k���Ƚb�i�G��0@!�-7��4�F��E-�����T�[�˫a��4��o!����q�v�D*)WJ����T;�9�a�Y�E	O,�د��dE�E��N��Q��z�LW�Gv���oa��@��V�oū�u��;\.�̏�uj����XI�"� ,��0D+9Ӡ�t_1%w#H����av�%�lH=������^��y \Ȳ��5�k���9P��d�C�h�6���}���K�go�O�d3T�o�Gw�/E�Q�.)d�������c0T��39������� mg�b~���[��\���f��v��>���w�P@��^�8��`QO,涨�;��2��2�/��ʞ����h��S�V�H7�� �7�^�(	(��ۊw:cƤ/�FWF�dS��8��=#���d�}�~�P��$e���{pk�J��K���G^�Q�(�v��w��V���j��<��{ 9��@تB���,%�$2��P�A�٨  <sM+�J���9
T���:􏡭������,�F&�|~�垽�)��s2�����XY��G�D9��۔w8�q��>�q@F�$�Z����F%|���W ��[;�m�߿�������یA���" �=��F'��&��Z�؉>�@��gs;;�������P]�#�/vZ���1��%{����e���]�~�/���Z���Gy�?�(�+*�!PkrV�h�g +�7߀3i|2�Nw���ʪ鲕$�9����{]�x�B���+~M�#'���#�VI�g�_�`�(���j �����zq��
�FɎ�l/��7�j���D��B�F)�^fl>g�Xm�M���o$����z�z@�$����SX$"����T�c,�*�W��^|(�<o/��u�sz	�u�q�Q>��=��Q�2��Y�v�^i�8�еQ�cs0���=�׼>9)ɍ��v_'E���`�ެ�73��`�i�f���6��L+>�F�ʔ�0D��G t����Ɛ���fۛѓ�Y=�dD��2���c�H�t��tN���!�oBK��9���pB%ҥ�:w�� �6X�lG{�<r-"����JW	�)���o��.�iL;�-�?��.���b/�g{���:��,3�p��`d�Ź�.:aZ�eY�G�NV���������?�_�R���_��H�Rd|���m"%�yt��6&P�p�U��	4�u�Xܕ������%ڮ�x!��n:��S����c���p7��
��y`!�?�Sr�@�Ec۽cMI�Ke�~� �q_~hBfL��d��Ukr�fH]ɚ����ݱ�;����
�3��](׽D��Qm��%M�=o&��c�&c���7r�P�ܦm��Ӿ����y��<9TǾ�xJ�9�q9� ��"w���m��,u(N�Q�1��f�W�܈	�i�>��'�]T��vCg	� =�$#
5�Pmӭ�@�_M�$�Cܦ�ЙU���6>�>���?f�/HvZB������3�-NE�˪u;^U�n1����F��t|��}Y��o���\�2i-<x�D��m+?Ǩs7>礙���*j����U�����Ҟ���)�Ε6�Z�տ��<���Y����0�r����a\2�m#T��$eg�rn��_���糅�-�[n�����.�⫊#�|��˥uBAE`�Fw_/��sxv����H��T�q�@��N��\�n�#	�&���xA-Nd��y�u;=���oc�~�k��s��j���II�}{����E�@�ߥ^��8�w���Dh�m����D]׹��|��2^	Ga��f�;�p�ׯ�؍_�c��ssX�n�^��-ty�+��6]�N��?�>7lZ���"�N"���v�0�y��|���K=Z�6|���ģ5��_���/�{���W����(R@���1�q�c>����!\�
�#""����3E��;���!�U4g���IkV�y��]M�w<�@���ӝ% -�$��O`����n/)���9kN̨���=ܫH�.�Y\L�.qd}O�<�����&�ʙG����z@�����z~d�@%w.K"rEbM�����}j��_�`ɯ9��mFy;�y)v^��(�;���#�%�L?�'Zr�D���R���Pzϼ�NVon/Di`�C�N���0�8{)cm�FEʷ�h���׏��C�'�8%>>E�(��o�/��o��
���a鸳�8��"�[���~Ծ�^�=y����MqR�� u�9����'�PMz��W��<�C�����4!��(�_��T����C%�Pp�x~��e������2�nn]|]�hQr���k��;��`)=k]��%�ˠ�c_%T�{H�#8����c��h�,�{�n��J���u�S�e���Ҷ���k��7T�cf�+κM�UI���OJ��C8�!�{�ۅ�V��ýh\��\�&�S��BhA�۱��A��0�g���o}�㱖�uU���㒶���J�M{8�Y4<V�\jiͭb	��ս��q�Z�������]�_Ih�uڕ�v[�ʎY�u������׋>�[�����+m���S#���bu�Ql�2�'}wP4QW�%�~�I���B����^0�HnY`��q�QG��!r��������/^�ψ�(��*O����v���B�ӿh͇�b
ri2O:���r
=��=��n�>fR�U�z:��N���
�
���m�G�T��u��ƂDt��Xe3b��ؒ������'p�Ԙ�Nh�-��w������g�;�3�6׋���V�CxH��_){�@�l�c�t8��U蛕��@D�vE�{�))��k������u�[�ؼ�U������s{GCn>N��'��x��%����%�z����kڛ*���c�R�1������6��/�m��Y�|�v��=J�Q�Te8�_c�É�Oޝ��a�4]��T�:7�I�b�|ѻ����9��Zb1�q�n�r�CC��6�팣�]~��K��5�KJ��u$����ys�V��-6o����|�#a,~&�� ��y�R�\��_����3�]_��[{��nE3YM�UU�V�m�/{����-��##"U�^婣�����R�n|����<|���NE���`c�i�ެR�a��G��&ؚ��}�ߏ�c������aƑ��V�������EjC1�l�(�.?�[�����vKv>�����
�����tq7�����I�����y~�R��n2͙���#j�0����@*�U�XT+�!B��/|���+�&vխ0��������{x/Ŝ��Zm9�|i��;E��|��4R
X=X��a�i���泉|�?ã�6ꖈ�H�>�RM�a�Б]�;�/
� ��uNwH����#b���USMϨ�$4�]�O�e7��iܘ�l���]T���`g���_%�/W�r
�w_���Չ��W;����L%�����X�_4����(���L��Z4��3\�VnG3&�8Ȧz��rf��l�)xhʻ�@9���= ����6;,����P�jo#VcѥA�Q9&̷�u'�
���e���@���
p���=ݽ�����H�f�$=�vQYR5#��q�>+g�:�<�d�Y���ҹ3�%����S�{ȊhL�㱜	h�G�Y����hN�0�o��X�a�4��@,��,�fٴ[��:w��3�Z"�#�]�W�#r�gD�#N���_SY\z�snL:�3��{(�V�������W�̘�%�T�f�s�bz�oˉ0�*� ��=lv������Kk�Z����8W�"E�K-/�E�2�6]Mo�wU-Ar��r�c1\Gf<�����A�6'��($@9D3������w�Y�M�T��|���:�]TO����f_Ķ+�~ֈ\�a�x`8���� 	-�[����*w�y�Χ�=�����=�WiN����i̫85ʷ���̼�@Bp�d)B#��y+�.�Hc��X~8�65��É^U�G�'����[n���^�-Vѐ�Z:P|Y���X�7	��m�;�T�l�d���8R�Q��? dϗQv0����X��x���;�]���t�{@4A����W�@�\6���Qj���B�]�сl�>�/�����J9���Z�(�i!n�铞�.8�s���J�y���L������f����0�`��f���u�k;��3��gJ1��xE����XG���3��
)�3�4~��z��@�ȋ�<��5��~���ķjc\�#M�?�W�d�c����(p|�!��޺�6䵪b�IR���G2'������[��eHr�Nz��l�^V�!њyU����ک'9��&K;n�h��Ќq	;���?��T��)oNӍ���m��=>��]6�B���|�yL�h�dG��8W���z~�m0��6�H\ӸK�j$�o��v}�!>�ⷖ�	S�UU_|v�.82�V�w,�l�Ġ	�Q����%�Vc_�ׯ��uǎ��-�<N@?����9���CqA����*�?S8�R?��6���:LQ(��zkh殰U���O>SuY&�����H�c��N�"|YD�8�h�fG�y�Ű��t�ј����gІ�1߂C���h@�9����jLo(ְ�m�Bl&C�rף��ߍ��^��i��3~Do�r;�CV��6CBI`�Vܾ��#qQ��Y�V,���~�:?���G���4l���4��X�$De�sig�#*��C���gj�JJ���ըL����%2�|~񞴔�����G�:+\`c��jS�6�-��V3��ʙ�c�׊&���s�.�t*�\
p��#׼7�k�����j��@]i7Jf�l���r�U�;@H�&�Up�V6(7��o����b��YT���l7����ф����U�7�a�A99tドF^wM�6��n1�j��r=C�B�����uX\�"�S�?��8r[fwl��}�%�h�KwM���u��E����pq'�wGt��R
�(���ҟ ܩ�]�����U��#A<�#(C(Dp���{ ���Ъ�1�����hV!WC���w�n��w����Iƴ��8�t��G�/2�8bL�A���s�naS���)��\��W�ӓ����6��9&Ƌe���=�XT���A[�n�.dZeQ�r����[ 9��U�ե�Z��v���`������:������C�h��3��`<ơ2�����BkI线��*�gxf��:��FR΀_K(މw�y.���e:E�,�M��:H�4���5��%���0���E�"ԥ~,*��*��W_#}pZ�K��9���yQc~26ί��SY�4�@�9�y?,
�OL��4�x?mZ�u<�Cxbq���(����MO�&�A�|��B 0q/&�4J�}2t�f��"��	[V�u�L�6��q����պ�q�mu�������Ol�#���Rw;�����c�m]���$pq?/�,:��aH	��6�ˋ���E���A��j���&�%tI��aC�:b_�;�d�ߎX!^�@����S�~�?6 !aWpM��]��K�/T�BH�+#rU8=�%����Jt]ĉ�Wڝ��};��x>;�5J���Q�͌\W��~�2��켛z<Ưnq��K����Lh^�������qf����|�&t9�����Y=����nZw�K�0��$J��e�s^r;%]w�B4�+h}�f,vï��u�
�Ȣ/k�taĸo���.��w���ds�1k�q(�Fy�Y��b2��rO�j��Z;xG�n��<�b�h�B�b�����l ə+��Q�n=⛠Y(�=������$�!%�n���TGY������(i��Gus'��&7�i�X#���������Ȟ�� Q��U����q��-d���9�J5�=�Ts���女���!���P����n,�(�r�h�q1<I� ��Yv␧qO��sA��Թ��Ht���k?ysN�愲����o��	���6��*�X*��w�gH���Q$�4�A!�@2&�����''�ӹE�バ}&�q�l$BnLMU���C5&+��0��h7�"*�������SB����'+��G׉�tC[�y�� ;j�v�$�Q�R{�ud����w�ܶ*�G�}�|�
�*(�qa��y�vPs�|�n��N���Q�5����p���`�������?77�e�0+��><��^S
?--��v=m�n��?��k� C �9�A� ��%<^�+j���@I|��m�
�俛d���f���tY߾p�y�fp�����pW��w@�\A��9���$��3k�4��hx���?�f��¸��̍E��}�]�ʨi�� ���u��<"�,���t�����h=�P��vcp*�n;�ʨ�[�Dα�M�o��U��zz5�E t#���=r�l�5D�y�H��v͹�i�c��z�0+����ku��s�zY׵���w>�7�~� v�W�섎�.e��#R�떧<��H2fPU�H(�|�S�f[�5���L�bϟYi�AÑ4D���	��$��#�rA��B�S!�n��J~G�R��w/�T$3�j
�a �Q~�ː�Օ�~�It��̒,��'�b�٬��D(dq��x�3���b�_l��/UHdH́$a^�'  	��T��%�������^�Xd����yZ�5<���=�'���F_}�u:�+��=��n�ayĆ�GX%}\�,���S���W7u������fch�o]7��!s}_��7�/8�d��Hы��2�*��@1j�F�n3{Go�I軠��7���z&k�6(���QO��t�ǐ�A��?C��@�Pb���	^�F�Bđ��Z=\.�����{?$3(�ϣ���S��Y�j�{z��a��'I[�ޟ�觙vy<9صh8mGX3�O�0<����!�x��d8O}��V#�;0�� Y�T,2��*�t_*s��FE{0W	������n:�OZ�ͱ���5���l��-K�	�Gk4��&`<�[lm��2�����4�{�d��q��Eo/�'�ÛK����E�=���UtW��{�(�nx�U�]g�N�%tԉ�O��ۙPq�W�%�
��Uŋ�<���?�3m���6�m}ϫZ^�dc��;K�H�h�hj��+\,dq8�
��J��ajW-s�.�-����_W�97H����L��{u+�^��&�U����kj�-�ߤ� :߹r���Ǫ���M_�e?"���>}�1gLV����/������a|�ƪ�q��V�דB�ׅ2� �d��'u}��Vө�S/fJ���a�@X�ze9�ͫ�wۿ �M��� �(C'�ـ����=����2ͱo�蝟dt{��l���h|�YyL��n�>�aq"��8���ú�O��V3��e��L�6��叙��,�b�s$(����o����-�xF!�:C9ǭ���@��x��M0<�	V��0�)j�S�� ���|A��Æ'�&�;�a
?��e9V��o��0�%���y �����S��*U��Fa�=c�Y>sQ�i1��SD>'�ڍf�H��C��4�[B;��@X	��^q�9'ݧ�$v�xqa�W����6+.DO?AX�����
��<�g*����E�����W��8A��s�?�޽��xUߪ��� �;�81ϑ�P��������6d���ަ:����(S�4@UFu��nCo=]������U����s�Zu=��v'�[M�!.#��,�f�CkϷ���71?��4I`��l���!��jE����(*�G������Go�]���q�q��k�3C���_-,��\���a�N:�"/ s��G�ho{� �M	��������]m'�aW���?��E}��˩�b���K�Y��	0"A�{�vL�XHLX���Q�#GUE%����\Z�+������D(��|AB�E��&�B.�(�Z�]6��lT����"N��+U�%�o��:I{��rCZL�i�\��6��z��+cvw�s_�Du����抖�g�����<�D�l����Co�~ztn�$�z٨6�^��q~��t��|�б������p���l�ǌ&��2����dk�֢d� 9Y�JV-��W��>R�}k��V�mݺe5��V����2r�m��� Y���e5�=�L��v�`1�Cu�N�( }3���m�6}�+�ݯ���)�1��5��
v������ڽʬ��PƗ4M	a�/j��ӯ�S��/Ӿ��KW��(o���o��]����.kNʸ6�?r�%�s��������d�7x��N6������䱼����#�?qC�)��
#}?߶�?�����S2m߮{z��27�rX�3rɇ�	G��������쏝�� �4I�6'�����斟�׭k��} �7�����@���WO��@�ok;�܎-2�3a9�U�J�(��$9X�?��7�p̨��yT��k`��8a>��D<�n ��^���f�fP��|�0�����r��s�A�'�m���B�a\��ԇ���P�	�� ��_$�9�����I�TB�k6����
N7��x|4�|a	�T����ϥv��z�R��<�����E���m��5�X>7��Y�AL���9�[��x�D��-z*�󖕻��}���4���[�%��������rp?�i�ҽ����KE?�2*��|CD�T��y�TT7C�������U$��gq[�i�;y|�Z_Х�X�qVE;�?�v�D˔��^,C*��tjz1J��<^����uc�Ei�Z���Yq�j� �U^YY��RtG;�w=W$ͧs�p�!x���8�d��L���Z�*�)�����o�9fК��~��i0:|-��O�;���[��%�v3x�4��˦�b�|'� )�P���Hdsx�{!Q�_���d�z��%��'�ɦ�%���� >����X"�k�uFT���̬��N���!��:t{6�&)+tq�D\�>|0������U,�$J��^�,3��iJ8"՘ncEķƱb �ʩ|��v�fY���{���t��%��ƶ�!e$�.p��0 c%��]�%wY��,��oC�-=WJ/"�z�	/�V�@�8'�==��x�o��M����|����@s�=��C��OZm}�Ï�7Q�+��o������?�p�PTd�|����_�2�?���vC�����#Fp��z$�=���]+k��>�O�``Í7�^�{� j��d�=��3V�!�|E/j��ۑ��,Ӊw�?i��4E�oޓ�8B�a�3��o��YH*	q��/A�C�����K^��/��ɫ;=��@|���a��A<B�~W%��Qj\P ����*�f�ml�؝l�ԩ6{��Գz��r�F���*�l�@=�;L�++[!W�ӿ�͟c�~>�f͞i�d�Ϝ9]�9Ӿ�r����3�2e�͙;�.Z�#3fδ��zʷ���M1�'ӛ2m�-��5v�O�\���MW�s��U��h_N���d�ĉ>
����'�|�;O���zL�*�(�Ue��[�**��[^���kI��/���@I�m���v��ǹ!_#���}Qf��fbtg��i>��f$�jF��@�Qv�3|/#jO<��Z�S��ϛc%V�����t��K.X����������T�6y�W6m�T��H���S��w߱���V(o:)�b���������{�4؎��O���\]"�o�8��/�'W@���0D'������޳%�	��.X8ߦM�"�,���q�>U�&)��w��g��Ï��P7Rèj� P��,�z	|�%jm�� F�����3g��Ӗ��e�#�Nw�]�i
�3�6��t��2v�ŗ}��i��+�(��TW�3k3}��_M'uR*Q��,���?�-�R���C��p�=�~��=��V�������^������_}�Ձ�{�Wŝ�ƣ�j(�g*�օ��Z"��)��3����aW^y�P��7ơϠ���\�~��ؾ��c��w��y�֧O;�gG�� �yD�a�W�p8,Ս7�l�?����3��!L�T����B���@��1����L�+)�d�_~�Ok�/�㢋.�[��W���.0}���~�
h,Qӣ���{�*Ӕ��V\ �X���K��A|�!�;츃=�����Իﳱ�a6w�l���z�}��&mhe��:���bTn��s?��۬Y�eD	H���|�b�$����`:#���e�-����O��(�2�C  ��SӝV�{2�0h})i0���ɷ�CxCgЭX.y��2MԳ6��2����ob:1�C�	'�C*a����BZ�w�u��N'�ĕ��UU���J;�3�sϱ�ee�T��o�n_L�����TU\�����jk����,ȬA*)��#L�
Sǖ��� B�: �3����Q��2e�G�$�DC�%�~�@$�w1͓���aĵ*_���:�YϞ�:�l��|5i����[VU�R�t�L�
�� c�����*�*�0��j%�����~���Q�8�'?��n����@�Fr�>1b����$��!M�6��1%��}��2�Uu�)y�qV�r����L+y��-3�Cå�zv���d'�p���<����W_��ȸ�֬��'��L0-�-��������#n�-�Q�:�O���t=:_�ߘf�1�>�<�C¦�V�lc�<�����8{�6m�-�)��u0���[�5T�%�>�Qu�����d@;���t\P~9.��D�ʰ�g�l�hvc�"������!6��x����| ��?��H6a4�|F7�p;ꈣ|����aS��ʘ<X2� �z�[F�
����$�+$�|�9~`驧�aw��7�� ş��(�=H-S�)}�o�OZ]��&�|[���&<���B�q�/-cq��m�'M��r�=���/���N�O����Os��[���W^ye��������_~ɺu�mE����0��
Q��o&D���UC�B�M7��N>�$����@�ʲ*KԈ�����ǎ:�(�ѿ馛��[o��L$д��;ֺt����~z���ϧUifۗ_|�k�ؚ�J�������,Tfj����aC��c_W[��^�k�0*������S�$Se֥k7�s����Cu#����{�����>
UP�A�C��v�<�S[ �~xu�V������n��Ͷ�N;;� �g���O�p�2Nv#����w0��GںN����{��,'g���ʴ9���y�]`?����۵kw�c4�� ���FtPzxγ(�h(�g|B���>��w1� �s�:k2h��_���xu�,�oG-|7�4*��,-�5�&�
����S#�O'��>�Į��~I.�\�/j��j����**W�>��������/~q�}1�_O3p`_5j����^�Jgzzg�*Z�L���m�܅��6[�����寷XEY��Y���^��Gٿ�{A�+� ��|壌U�!Nn�@��Qq��Z����o�tdؗ_N��?�~�#�P��[��	���@^��]w]ׅE�Y��2?��{�v��g�a�n]:����~��~ڙ2|��G?>�n��Oֽ+�H��$I;�Q60��"�[v�\�#'� nQQ��2��������,Y�āKW�x������ӽ=f��I�2�??N`�5�)/g�� �g 6t�
�� F'�|������|�M�����wߗ��ǌ��*� 9�)i+���n��j�^�k��Jq� �ǪsX�f;���z�A�<�`yi����zV��A@��������9�m����e��4"Y'��"����05�]� $��	����6<c[��|ʸ�Q�l��n���-�1�U��K�FՁԇ��L�f�ӰaC}���q��(ӌ3}Z��o!�����$�K�B;��Sm��v4��ʓ:��t�����(}�8�Z�֛�Ĳ	�]��CӚ�%�<�i��m���Ϛ�L}�Jm�p��D�M�:������7�tK�޽+����ZLߟ�ӷ��ʪ�g�{�G��Ϳ�w�����O[��jL�zC��V�2��BG�@����g�*+*S:��jcWz���g[n��u*�f�+J�Ѥ�[�|�=��O�q��@��f�mm�����f�j�+i���6l�H�[c�-�a[�C�B `�6��q�=����;o[a�0����w��6c��7z];��C|�"���W��aj�6��1��1������[nu�}��I;S�_���ox�h0��+�=�ܥ2�b�_w�oT�+g���SqG{��w���}*�Ʌ,y�v������>��3�g���~ݺv��k�V�,wЈ��<i%����.6B���� <\�3�Ix���� �q����Ȧ�!d�3��?�gz"c�w8�&viƐ�W���<�iUer:��o�?=��D���T5[�eF@1�I��ǙL���>1���~�l�x**�񯶓N:��>��B��/ى'��#�o0�6�h��~�#��K��c�=�J�s�-��#�=�pj}�wv���xݻ�q����>ա�غu�fm��}9i�����#C��{��l��(�y�P�w�^�i�QG����Gv'(���O��'�|���d�M�5����;�m�Ŗ~(4��<����{P=Pf���b��_Xan����ة'��8�أ�뮵.�;����J. $���Ju��׷O_߱�uK�������VV.�)�0��U�e�uFY��ݰ�b�ͽ��Q  :�2���X�2 �p�k�OaD'�t�����t��|p����Lq{�駼n`|���8���{���l��v�#�<ºu�꣺L�{������2�|�~�p��\W>��S�ٴ�S}�Gy�z��r���=�P{��7lР���Nc�~e
ӑG��;�1eq���>����6�)�Ç�(P���An�n]0����ZP�:33[��eJ@(;��0*�sИ���Ξ;��κ�0rő춷�����o�co����$�w����_~��V<a�D�<�K;�³�7�^.>�Tר|�f��w�<�� yC]�\��#�FZ�r�o�P����K�<�:�g���}_�i��ք^��BH �u����s�̮9ꨣO��k�S9�i���9�N?8�u�م26UE4V�vє)S�H��GL���r�k�x�o�.���t�T�ormU�<�O��0��G�e$ *���\�~�v�o�٢���+!��P�]�@@�o��ڄ��{:P����7f��b�(��_zp�A�c���m�	^yc�@���p���oF��C6��������v҉'�!d�;�xkl�.%]l����C>DF�&�馛�{�a����מ2�����fw�y�m�ц��v��T�������2�`@��j�)S���a犞��2�޽�m���v���!㴧�ְ����+�;���@���m��Ʒ�挖Ν�}���*������YU���(��	@Y0n"E}���ót�ߡ��(
#H,�˖/���v�e'���b;ӵ�'Cz�@�0�p��ʁ�C��-��\@t��`7}�I�[W�?����Qb]�[����1b�O�am�֒kw���{sd�*��Κ�GLwbD�k������5ε�w��j�#]舃!��+M��Hr7�_/��g=ZBF' ��e�M�*ې�f5��^cl��f��������3��SO�S�6X�>�ddn~𱕗UZaA+�˵��֦O�i˖����F�޵��h�{���b=_a��56�� 罪��fΘ�� ���YO��ڥ�J:u�a�:�6��xϝ;OF�t�?o���96u�4�U�����fΜe�f��m�?��}ﴨ�X��f�-��uF���$�ز%K����}:Χ2mj���M7��i?~�=��d�V�v;ni�ﶫ�6��)��oxY��a뭷���6X��F��V+��v��O��׆�2�Kr���!~l]���[+O��\��>�׳G/�T��GH:[�GFFJ:[AQ��Q�"p��y{�|b[mt`���i�>�Q����f͚�<*S~}�#,t�Pw�uW;YuN���������)ӽn+((�9��W��y��n�+KW��A��������=��g����:�뷉*���/𩶋-���g�Y��]l���f�}d� ������7�d4 �9�u�{����FɃ�:��0���d���j0�*��*;u55V��k��М9r��S-s�sm�����m��}��������u����H�����Qƅ�ۤI�B�|3տ���2�Y~E �i�]U&c��P�hwT'EK�L�cޭ�<�'�V,é�C�[(��@<׽I�L�.�5�O�m��U=Ku�)��߶�WLS���xh�T�V�+ZUX���c�΍���E]
������f�m�i����ꪫ�;����iO;}'4sƬ.����Q*T�<��3]Xd����a�BT�P�
į���fg(��)�WkR�I�ؚ ��J��upe���~�kz蹝<e��'۽v�|@����1B9$1[F�3a1����,'������~�=����K=�( ��
��V �Ԡ(��+ܐ����{�.�Wa��X�8��d�
�A�����E�vo�R&�����t:w����#�8J�Ǿ	E4��<Xc�$A�z��V��`�c�WHVǟt��z�I>5���7q!z�I_~�kO؞��_8��0}����.Z��?��]p�y�>U�N/|�;���oK�;��� �Ţ�ehf����ƌmU2��b�B���Ե�)_ &O�x�͖A������:�{z���,`��dd9Y�`�-��Ȕ�:��Ry�8e�}w���+��^|ɺ��3=����0�;A���'���2;�G?��O;�e˂w���t��^z�~��_�:��Hgl�WG��2�*�5��㎲c�=Veb�}���v�'x����+����`�k�q�V�]҈7P�}5e�o�A��hfM��LgcĖ�'���FM	��@�z�+]Q�q�W
\����mg�q��k!N�������r�M��m�}��'�$���{O����
r/�������v�	Ǫ,v�;��N=�4�Uv�E��%�\&������3;��#l���6r�P�a����H��W_R�H7r��C� [��6l�d�O:��?��=OIg�g�Dm]���(�2�W�I����$�{B�e�N
��2���6t��i̘������Fm��Y/X  z�U��8���1c6��?>���J�T�j<x�u+	#H��}.'���?�P��� ��T�!k�2�^a
"�Gl6�;OW"L!��3��B���5c���e>JM}��.�t��[�BuQy�˔]6��B'���-���Krl4�v��m��F�e�oq���G(�=�.��/�����Ϯ�g�q����[mؐa.�*�ј/�+�٢���҅��2�6���0S���ih�X�R�<�쬎"��D��S�=^��(�ٕ��,����VE���+���T����D�"MJ�B[M�,���Ǚ�����5�&�h����G��2:�ē
�ϟ����?���I��T�ѱ��ĵUY��~���;|}
߶P��UQj�k�M:���������e�T�.uG�S?�Ã�c�F�
�a1P���@d�r�Qe�S�X�LCMc�񇁊���)������Bc�Y@-;�񌆔< m��&~��'�|f���������0ݒF�) l���������o��~�Y�^�L|3��0&}�����j�C����;��
�1:q�/���N�{�6��;u�l��E���ݛ���0<�����/�"�I�x�駞�Q%v�����jТ��V�O�|㢌q� !F�F������v�� ���86�`W>��)Ӧ�t2FF�xNO|gw]��%�;[7��߀#�[�	�L�� � ��n����$l���6L���1X!�m��Y��
8�Ѻ���J:��^Sc�!S҂�w�aG[�����-����������ys�!�(�(�T�Y��.QW�l��7���l�r{���Hʽ�)N�t������c D� 7���U�y�y[���<Yn�
�e��,�F�,9'g�`� |"#�b0�~��d�M6�M�b�
�z?�rɺd۫W_�K�{���|$��|��� 3��F�K/:�{�l�+͊ٶ�vK�~�ҝc�,��c7���9F�:ۈ�#����\0��Gx� � ����z�m$�����E� ���|�^{�5/�o����}��������^b=w�\�'�9Kl���"l#Ύx�mʔi�6�l�qA+V�z\��#��}�E��>R<�>���sy��rP5�u�ܹ��G󑳑�eV�:�ؖ��������)j�!���YB� x���$������k*o��f��������>��=��3����^y��8��٤I�m��/t��}S��ԩ3}4q�@�� �;��7�Ȯ��J�G9d�?��^}�U���l��˖/�]vk;l������ў{�_��bI�7��R(Sa�$��@��цU�5��k�B�1�~Z��.���t/-�;�g��{t#�[`���!iu�gH6�����C��:\�9W>�o��O���[���S;@Z���O)P���*�� H� А���h�Bo����hU���֠�k��6���E���U�w��h���g��2'~�wt���'2
��.�%[벻��F������'�|�^x�#/ F Q�#�\��C�O���wFn��9�1 x�a��ƛ�;o�m��w���b�`�ϤI��7c�ͷ޴	_L��L���K˖��h��:��s@���YVv�7>1_|ʡ�Ѝ�����ȉ�Il�{��'[^A8���3�x�M{�w��>�����!�!F��������VKu��ēO�A�1�d�T�Y48"��ߑ��hty^ԡ��m������g�9�T+��2���(P����������]z��Ѓ
���
��n(#;�j�{��3x�7[i��λ|q:���!`q��a�};�e�e>Ň���*�}�C=b��z��eE�l�^V^f]�u���;�v�e�=g���pH0=������o@��/^�-^qŕ��'<�L�D��5� B>���|u˴,v\c��Fm�ӯf͚���T�T
,wH*���W�U���=� dN�����f4�X�FX(O��Vz�!e#�~�PxaK초���)# Lg�0�X�����R�)#��G X�6� �b�.��m�Ֆ���@���@.Q_m�Ǭg;��٧�͜=�{�Q��2�*޺t����H_���'��ݺx�H`�1�I� #����&���# ���A�@�F�A�}-Uq�^NH{��aMSF�'�E���r�4z�7'�p��;�A#�?ȄM0�T���p��B�yI�DvW<l��YRS�}L �t��5�>� ˗�BL�{���R#Y1��O��7��,���#�D��): x�Q��C^���hG���Or̒N��%:\�l���Io� ��j��:2t�3�� �N�:E���./--�����pG�P�-Z��v�c�v�<~v�|���T�|���DS�
<��P_韨Q?�;=W������:�/y�t�w�'/r�㓀�8�Q�5��5�
um��5u�n��T�3�jyK��- �$�N�U���S��|2Tv�p��K7�x�_��I����u�ԊT�ds5U�����h 1(��rIw�Wza��߯�K'��O�wEk���)L���ha%������z�m͘:y���N�NÎ��E������V�k����y����`�O$�#���'/ᙆ���oL� �t�L�b�h�ð�S�h�1~h�٪�
~X��{�"xz�_|�E{��w<z�1N�ǵ���\�U�҅�.%�AF��hGq�����/�/���=�\��o~g�]���م^h��~�e\����h�2_����|�i��b��e�1ʅt�����5����gt0Г�'�
$!_�-�:5��A���;lƴ�n�c@FXb��8�H����\��{�{�H�=���[oq��4[ܸ��AH�����@Ԕ)_'�ӻ�jjL��Q6{�B�g�@�:͠#�PϘ��("��(�Ì��#�cmiǨ$mQ���IwP|�
�8���FU����N��(�Z����(�I|����9e���J�>e@�`�"7�w�u�⡷��������O�B��`;�gc�k���-����n��6��g�I TEE�O�b�4�l��������"�������(�$=��)��$Q��0BRYU�y�A���F�'\�0���F�gL�%����c'L���&H�
l�}�W8��̞=�e7z���<��O��wLI�=:X���q�{� �x���qC�Ǝ���P� "[���3��B��(3��|� R��7Գ���AW�#�ȓ��A�˙s ?�?F��H:d�p�L��Jèu׳�~v�{�q���.��T7.]��u��Q,�Ś���B�g�򥃃j:OD� F�#����:�>�X�'p��!Y��0���5�D� �n�F�Q$d�����;>��\�㞑O���_~X�G��ۣ�ԟ��=�=�|����c��=�F��Mx�]��������'~��oIw����E�Ku�v�g�+Lqe4:���F�Pq�����Q���5��UIԄ�-T�C�H-�m���-k��	^V�R+��~8j���q��c2��(c c�y�]���1l�٦>'��K�
��
��~��o�SY��r^F��E2�1��a��u��b~�nĢ�Yl�h:�{�M�H�#�_�#nn������f��n��
�m[��
j~�?��|G��d���_~!v���>lw���޷�ez S���� ia*�g#1&��5��7��t�R��EJ���3��a�H0�0���iMM/�C��d?B`����cLD����:d�0�r#��������1��-�б�ߗ�, �� ��8�@�u�?�7z%3�r}� �g�K��I��	Á��.�o"��1�aa�0e������uY�����E.���� �t�'F1 	0�$M��h[�e4k��c��~��|+�~خ��J�|��W�)�������b�f�p�RȎP����
����JW�����X�ƹC 6E!m�5�A\�rc�xyF�y��:�:/ǒA��aĔ��5�9�<�z���:�nw���y�.p��_��w�Ġ��8��ᶿ�!p��]ݟ8m�ɦ��3��C?d�<���p|��^={+O�|������'dQ�4��KG� ś-٬4���?�'u	|�v��������)��7 Rj i$��8�?\�����od@�Ȅ�x $��S����1�ϴ;F�ؠ䮻�^|���N��i��v�-���v��念v���7��.q�KHc���;@ l��1;3���-k�"�B��@��ư�8�!s$�PN�wN8��6��q:�&��,��;�����{��
1��\�e�y~�c�\O輻}ͩ� �ض!���U���ᾄ˻�!B��o~��\#�%��9a��?8�il�����	��Gيe��"��<���
o�E� j�-];��4����ۯO���j��be�5�bALu�Mj+�t���)v8�gn 0pT���=��kB/'�amM�I�c�S�X��s�6�0H0���]��5�'�aLj�#z��`ô�E�{?�ت�8ᗩ9L�����H��o��Pi�F���ք��8ܖ)h�:������j�m$�b7�ص����Bq�iA�y����Q��I��z�:�:�pU�G���3݁��'�w*�b9C��Ć�1ȹo���E�Ɵ!;�k�P�ؠ3���Y�CT��^0|D��B@7�`�ӷ��T�R<8�2�Y��1���I+a�D>�Sr�PRI:�!���Z�3���!�1~�� ����(g�G��w�!��c�a����Hi��>}z�_Lw=���{FS�sF*T �}�����3��02Q���<gHWk��e8ؤ3�ݥ�]#�)�"$ Ж�E:�7��[�NF�j�-L�Do��uF\����;��`$��@v�_�T���; ��˸'}Ld= ��2J4v�Nv�	'��HW����z��dô3�it�0�٣�u���7x���
H0:��!�6�6 �`��G��IO*��lW�$�/�F�?:I��!L� |t5�Ȇ�E&ć��gZ%�!�3��,F��ϹD;츃o���{��?>��q�=Q/:k��t�͞��u�xq��I��Ag5���& �B��<�������ors
j��Qa�	�e(^���>�G)Ic�ȍ��z�ox�gܻl�\:��B�Ǩ!�|��y�1���e�N6�OҎ,^���;�A�,d�B�ԃ�8���m:C�b��^�	݇g���=��M�>k�gj�hK�z͆GL�� �X>�+(��p�A��b�
z*E������J�D>y���y���6��i��v���*��	/��G%�� A�Ku��D�t[nm���K�{�+lF�Sg�Fj��0��
�J����ʞ��J�
�]� UL��B�Bެ����cނE��ゑ����� W�nQhՠ����=��#�'6�P0 ��l�#����;�_�re��N���i����f�{�c~�T���4����D���Bȏ��s�VG�����"������k�Lʀkz���{6�@f�d!_�qm&?�CCq�$����c�Q�S�040̘>� #�`b��C��xQM�+��F�OѓC!��t[�{�B���(WA��	��h������$����3~)o<�F�O<)c�U��g;�Ȕ�_z����[=�<�7����4T����'�f�-����=��r���� t�� v֓ .��@�$��a��6��.�A���$ �R�EgcxA��,[�B���e��� ��X�EBG:I^[m�����+
��#���T_t��v�ig؇}��8�b��f����H+S�q��L��Z�et�i��n��L�u���G]��2(�+�[�cP��Xgr�t�ty�7�#��A� �G}��B����?�� E/����{�~6��/m�����v����?��t���ފ7���"�X>�5ç�!�+ 2��`���!��α���}vf�u��݊;�P�K�sKt��
�:��p�W+r�:4p�y���G��h�`�/׶Y�2f����>��Mb8���ZF"�T�={X�.]��>m��J��fĈ�6h��0*+�˚VF<yΆ6�r�-3X��li��L��ӦN��T��9]ȝ��9sfY��⡓�6�����Y3gxہ�P��#(c1�����8 ���P�%�	��:Ĉ�ң*;�e���#
5t;�U�®�jm
�匂~y���}x﯒O�?��չ�B*[S2�.�t�N�_X8��������,R��b��l0"0x�1�bg.�D�D%]_�pC���ʚ-��/�A0��t�U�'"<�_�p�͜5��>��G�X0Δ��3jC���zv���v���,X�,��+ғڐ����wЗ��΍=op�|��,D�2��y*����n���b�E��^B�ö�|�?g�Ĵ�f٬����ז~�4���k��#�Ң4�Af���ȑorGȏ+�=4ΑZ5��6J0��#6�d�[!ru���]g�Xf����E�e�5,�q���.Hcw�	��6*dΨ��24I7I[Lc�۷%�B:I##���#!L��
q��_+^1��X�5�B��F�#h�lr ?~��8�����H(��0j�Ƣ�#~�L�T0�
>	��)���5�A.Q6~�ʪ���� �P ��9e *�{P��1�h TUQ���r�8I����<ݤa�Rs�+���ŕ4�QO;t��出��	�L�bo������i�p���U���]�ܝ�'��o�a�� ����{���ys=L�R���J#�&}��`<��aZ&e�$���'�@d ��=��s���.��U��y��R�?�1���t�x���[��7Qw��n��f�ӟ�#������.�s�?�-�nݻZa�B�8�r�*B9,�_҇#|t����vء>j���
%��6i	���Q4ڇ�*c<C�s���,_^��j����%�2��9�;���`ͨ ����'�" %@�z*ԇ��#'�R��{t|���,*6Ĺ��;m�]vVg�4�i�/t����G{�~�_XQ�b;����?j�=��o�δ��_�>{�����K.�Q��w��|�A���{m��w��K�T���_}�|(�K.�Dq?.��DBz?��[w�]w��
������bw�y�]{ݵ���z�0R�, H�GG!m�ZX(����]'�f��m� 6I�
���mYЃ�68/T	ɼ�����v������V�*�L5�C���	S��H7����]�^gS��L��2�}����9Γ#��|��AZ�[J�gU���P�a��ѐp��xv�iq�OTQ�1w��G�g�T�"^b�.��U�yE�X�h�j�
r-�I���s�8�ÕF� ��0�L���T�WP�'��e˰�e�8�5�2�,K����<���F��lV0}�4�X���=�L�ԩD�B�=�[4�2�dL0mE�n6�Ab�ӻ�l�/��C���I�*m�ѱ�d�Ja4�]��Б�'2�$���|K� �<.��&;�2���
�X�c�`����{�0�9��%��H3�Nw�<Dǳt���o���Oz�g-�!~F�}Ue�����#���8�w��'�d�0��>�y�Pb�A9�+Y5�h��}�W�W���+�j��c��7�w�Y���/U�	��}l����e�(.��B���Qr⎠,U���"-�"�&:�A��+��eS.�� n�~d(n6�@LU�9���UV��TF`��O�ϡs����|��E��n@�,-��eu�X�C.������^h�]v�ŧ�]/C�-��a���� g̗L���"��2DU��K����la�����\z�TTU����{�ceie3�_�x���VXn��W�ŋ�������NXm��LE�x�Q���־�^eF�˔���-�o�cT�xf�
cK�]��s�'��Ie��
|ʰ�ٯ.�X2Ȳ�n�U�z�˃+�S�s�	#�w �g���ױ!CFH���s�w�2�c�HKY�8�5�H��� �,u��S��g9�u,GQw�b��at�����;�-S�:D\p��>��=��>�;�8���,7�W�HcU_F��w����W��R���m@���4�T��~k�3��q�vַ_O[�t�>��Uz�)_0FJ�5��f͙f_M�B��n6pp7�	�VP�h�K���韫N_�:p� �b�i�ٹsXE�����i��,�e��.��.�5*���R��m��y�����W��>j�2h�m��z���ΰC;@�bw�O�	�~�mm�-6V������׆�o���al��F�n�l�����r�l�F9�<x���������޻�UW]a�캓��r�٫������_�o;ﴭ��^ֽG>b=��ګ��ӎ�����~�����c~bGq��}��v��lGy�¨���u���icS�����l�.Xj�Ǭc{��7z�ʌ�Ty�:.����6�u&��}�q����t-����hխd;�`�BU��AA�� z�K��k;���Q�Su��	��ƙN�g�ɒ��#���1{8!o\�'&��h���e4+LF|ƪ��|y~���Ĝ�j�d=\���-��Ƌ��(d�w>�#n�ڣo�+������VP�9��>>�����QC��e�)�ũ{���|Ooz�%qa�`��V	c����Ȃt0���Bx!n�|�"��;�#�7W��A�D��_�L<�� �B>z~�p.���m�W_�C��x���򀸆0���'��=㊼�$��Æڶ�l+�Uٌ�=|K� *�gD�u/��I����}���=���eL7b����]���.F
p�F�I/S<Y3(i�y��Lz�g4���{tݷV.*�����&����o��XY����Yg��F3���]��O�Qx>%9����0էw7\��R	`������K�ҙ�הO��r`�(��G؎�m�k=���9�����	�z�<FN��e���2J���^1jG]y{챾A�9�c�=���8�tR�����^�zڠA��W�|[y�AG/9|�<�/S��b�"�DZX��SG����u� \�E9�.��Y�#��80�;t�G�����l�����?��G}čyFP�.HGӿ�5��,OKyY�����V��w���:xñ�
<H�v���y�γ!��Q4���Ug4���y��C|z|�QGI'�MO=��=�����'����f??���
?R���~���l�6���e��0jrɯ/�k������ �$lmN]M��;�z�J�G��6:�8���߶�Sg��6r� ��b��]��W��������:�	C�olq��'��'gG}�s��>���I�}���4@F�ٹ1���6\��>�ē��_.��o�R�QAa���cm�݈�l�����?��^~�V�-֓F0��]v��v�a���e�	f"̙=��2M�2��^!��mC��y @!�P(*�=7֗�K�3�"�(���a��R;@Z�H�y���*Tn�Q�(`�����N�&�t�J4b�C
��W*X�h����G#ȕw�q#@�g��{�J�'�S:/�6F��==����cD����hLS�~��"n��`,�̍���c��{�c��Ǖ�URD��W�`db�`���C�8`č�#Lb������}�D\��W�F��y��.K�)� W��&�κ�}+e�U_o�h�K��-��ť�"�?��?�D�B�o���6`� {����y�1ސ�'�~�����`�oS�:_{č����_	=r��<#�q����� �P!�1�I:��%���n`� l2�?��9�[��Ȇlg҉'����n��ü��}3�#l@�1��t�2��I��Ec^�e02m6�JLO$��2��v$�[�ZԵ{W5�H���q�WT���)��QV��Q5�=v΃��a7�,O~#��(6"@ج����f����o���8(�ukg�y���LC�|���ޑq� �@b���z����(��#�K�.q����b]�w��}��0��VI9�e!�e�
q��;�ߩ��8���_2�u��Z��_^bO>�m�yqlX���۶�mc�����y�M���s��7?.�-�2�|�2/k�q�p����H��m��6u�,ũ:��������^�S�:1H,{X��ǟ`�\s�m���:�l���l�M֗>oj�s�]~��l�H�L��l���;®��r��R<�}d��3ϱs�:�~��s�c���J�d����'�n6�x啗��ϷO?��F�,^f�+�����u� ha!�r��	>��{�����C��=w��� Vք�_�7��� i�m�������
��e������Fn��Un��F;��#��~f�]�-Z�������9� ?bb�ܙJ�
����;X�`ɍ�I�6���".t���m;�ӷ�֭B;��t�B5�}UY��ېB42�R��VM�'�!?*�����	�V5����=��Õ�=.��ѡW*N�H��H� +T��vV�#��Ϲ�q!�XS���E�bi�#,��7z�7�F�~�b�����@"�����Ϸ-a�5+2�}$)SqaH5��K2��e26������∏0�Q�����h8�	�1������Ӆ��tҚRj�ȍ{�	�P ��b䈩(���sҽ�Nc���Hyܞy�I����Cۯ�k�&�T9B>��E���L�����|�D�[��������2p�ӟ�!��;o��}����SD�7�9�t�M��ӷ���v��RP� ��o�� ��n�}�ܠ��#���������G]��o�Gw1�8��Gup�a��!����fw�y��@�%��8�"�����'F��= �9��\� O�N��5�ގ����ʐ�(�y��� ��qҗ_�������]ب'�C���>!#�)K��7����wЈLO;�4�������]���o?߹�{��#vu#<·��O�<�Oȅ��8�G�/�����|�M��h!�M�a���$�Q~��5�������;��w�+~�yO�Q7�}���7.�{�W����n��#���d����۞���v����z��V[�N������'�?�H���:t)��a��Ȅu=� 쥲w�G�.��n�&M����
{≧z��
55�ʮ��5a�(����8H�C��&L��z�Q����}�)��م]$�.���ϖ���v�e��~�<�����*".d����:�!3�����Z�i8�I�|��w�+����p�q�2i�靼�ݷ��6���!�|�i�7ѫ8RC^ѹȈ2���/S�KX��lp�gu
�)r<�g�=���ܧH���ټ9�얿�n������֏unŝ��)���<��ϕ�`��k���;R�T��u�δ-�҈��%A��.q5If1y��?@� i-#�,5h�8d�@P�Z��`���"�b��Qy}bD!=��R�����j��T��S]$�1����[�=�4� jW�*Y�J-�t@4����D4B��ix�B�o���k�k�P��=�&�س��!,�c��ǣ�|���(ӆxN\�� ��f�#��^ �'���L�~Әb�W�R��3IӤ��5'��K�L&�;$�1|���&4E�Ƹ��˞n��zjDK>����"�W4�p������x� Z�1�t�)M]:۰�����}lؐ���:�����}jiA��	G�y��&ybd*����_|as� ���7�p[���`E�ؠ��C0 YsvϺ��lH��x���g|��z
�g�l@$:���?ҁ!�Ț4bTc�3�d#��˝���;�w
�+�w�a���o��U�^)�/��Xd��1���~��}:;%R�[������O��0���	e�o�?��=��ȝtWVV4�kvx#�!J�`�\c�-���6e�t�3g����Ǻ$���#S�9��n�J�uT��{�½��{v�%��������u���Lw:����O�����1�0b3�H�G�� #	Ȃ�\gϞ��+s#�86�q��G����P>�6ᢨ�[�ǃ`�W*Q���w��	���y���m���'�O�/�y�<�"�Y��[n���>�l�����#����TY�k����0v�C����͖�Ȑ�F��&�g�?�d�[�b��ٳg��
��?Rng��,�Zgٖ����ގ�z1:6�8p�?�:u�'p{�QG���i<��(>�`��2�G�z�!7򫥏�^{�b�^v�|�l�vP��:Rt��3U�N�h҂����>�A�	�3�6��B�\{� �JG��h#�i^g$Ajl��'35�s�.6b�;��S�?�h�_x������8�/6'yD��0J؂E�|
ᗓ&y��Gα���)R7E�YI�ʫ*�c��͟�@�/���.��%֯Oo˕>������>�3�+�I�}Dܷ���+j�"C'�;1�p�C����w�@;}����2R!c��|zvih.�� .�������I�����OZ]�֔���B���nQ��.�
�l�t1���#i���$?/�Z�[x��ק�ɏ�$~t���6D�4�ć#�<��aPaX`d0��+q`��>|Z��c�`�ѠbI��=�
�yUD��<���wK�q�g��<�ƕ�1
	��"G�aa:<�u(�c��=@��R�=���E2�����\�,�(�_�3Ҩ�68��CI�a ?*���e`M�1�f̚me`��/�q
�#�8����ɰ�Ѣ���-F�l�c�u[ٹy6j�(7ğ{�y_'k��{�=j���^!7FF � �.�h�C����$�����re�x�LN�2��>~ �k�c�Ч�~�ϑ��5��sf��m��GW�9v$ /���C��#.��{��{�
z�J��=��0�%��+UV�AY�S��k�8_*��9�ɼ�O�����Զ}������|�͕O+}G�g�}����A `S�*}3�O6QV���)u� T�ca�����͐NR��/ �D:H��O?m>��_ZtԐ&��0"�2�"���]�Z��߳�3��x�D,h���#�$�Q��r Q΂| "_p����C�	yH؀$��� Ϻ�7�7k�@N����vƙg٫�~����iS쭷��m�	�os��N}�G�#`W���N����f�Ѹ����{��_��9[�?�;Ж-����5l]6���у�¨��%�m��y���l�!��aD���J8�e[q��0�~��#���o���:��/��h{H�wf%ˑn�>Z��\�r6v�.��F�Z��,)�&O�g�{�x�{���V�sP���F��J����m��Vv�W�Yg��zx����_�?��=�#]��/i'�p�x�<��Iu�kQW ��y|K�6&[mm^��&��0�c����δ;	�����G�ǟ|����s³�����Eȅ(�����F�"O��k��(
�i\%]k~�Nk?�����@d���ZϤ�(`PK���1���%�G8DL/�g�1�
����1�Fߧ��� �q��"Ǡ���ݫ��q##��"�p^JxF�L� ��x���p8&=c6�A���t�8�=F4=�L+��w�=��l* \�*E]j+Q�P�ӌq�˒.%ֽ[w�-0.!���0��{h���sk��rK_'AǴ0�E�2^��ABV�E=l+��Zv���9�W�<�r����� �I�7�zSF�iv���������t���M7���A�jl����|z�O���zǳ�v�w�������#�ɑa�T�����#g�אǄ��^{Y�>�]��C��{E⿿I>kLI��'����3Ҁ�Q_�7Ωa�G�@���9AO�sdGYAQ>�:��IϽ,&�nי��� �0�1�yu�{G�+e@��"M�8�O�e��⨈�m��0���3y�W��/�y;�<t�03f� �{���[m��Hgs x"�8�( �A͝�q��Ѷ��z��v�it���h��3L��h���kݱ�5�C���E]�S���sO/��E�L����!�=nv-����K~���Oܯ烏�^g�H�.�AR]\&�J���~����| �Po2@��G��k�������A�W
�4 �r����s�˓p9��k�n�3�3�4s�L�"���Dꁁٌ���O?��G:�3u�>c�m���v�I���?�����������ia�!v@�����i��Qv�9gک��nW^y�v��JoGW^Qjεj+N:�$���?G��X�,�B�(���^�Ļ*�<����֭k��T��z�9;����׿���������^��9*k̔��kP�¦O�iK��Z�����^:Т^PN�t�?w����;��g�5�ob���4���7�0��*�)ԡ|K�
����v�i�����:�L�@�l�V��E�!��(����B���e�N��R��ZAjD2d�4Q���)XјK-��M�>��7(T�4��:�:�ӨӀb�Y��⋉z���0q����J���q(�E���a�q n��;�J���)��Knx����d�i�d�R���9�Şi �7Ԋ��ㆸh}�-���Х�"E�� ��`E8���ߧ<a ��Yb���H4fP�T��S�}hU:�򕟘�M1-�"��T��C6
_W�������o۸O?q���l����k�ۋ�FH�E�A�-<E�_�!���7��3�r�7�m��m��f��쯾���d��x�S��À�[��}m������w0D.K��������(S���v���fx���-1�H/�qvɗ_~)cs��D�#��0�/���o�\FP ԀF=S`y6d�L�b��!����޾5: ���c�ڀ�h�G䅃����(?�b�5:<��T�:�ҡ��H�u`���}�@FXH��\�K/�����[J�pr?��/��]p���ut�/���g�9�1�4~<�?��:�P��ؘ�s���������?�?��_{q뭷�{6i����k�X�Ĉ��]�.����o~�k�x��)����������nk}���|����mĨ!����8p�3�T���= �H��Ʋ�H��� W@'Ŀ�V[y���~���R1��<f�2�n�l%L:�_f̘�H����(ڍ7�dw�~�=����c���������A>th ����eǮw��=��#~~#>8x>l��J�]�����L�?���[<���o�3|F����_����:w�SO9Ѯ��v�	'���֓��5��{FB��اEfK~�U���W_ظ	�l��EA�� .�S�D������/t��6������{ᅗm�<63Yh�-�A��WT�I����������o�����)ҫ�\�X��hb
u�9����ٹ�Y@b�:b�G�"��P��

s�GϮ
#C��� ��SX������X�#�z�t�
`=��ԧ���%�Ӷ��qĈ|�Oʿ��v��Ժfk��d<&�U�d���Pq�pQ�|���
S�8o���};J-�~M�G�r?$E^#!���}X����	Sh 	Y�K���Vr���~3�	#���9�U>��X�O���QA����sƉ���L��O�T����֩�$Lz���I������)-8z��M�i�apGc�4&~1T�*� �t1�{\��0��R�'?����ȌF/�b�O�>Í'�#s�'O��Fw�}���/�+��jO<�����{�'����F=D�Ԝ?mP|�*?�ϣ�@��.�.ȳ?I�)6z�9k%<kpR"p����H�Ț�8�@�]���NA�@�~�;0�ԧlb��koʨ���pp�l�Ap���^{�'#\��;�s~^^�O�"��ϑi��o˭	�����M�tOaWV�Ƞ["�o�-|YG0w�|��"�ַV�g̰�>e�2�`��e��z�7�x#��mݯ+��[��1c������H�������a�Ȗ2�De�ʈ�u�s$�9s��]��a2���7߲7�/^��H#��tJ��D٤��羖!��[��m�y���H���4-F��,P0|�0鐌��]F�="��;��`��f7��;܎9�g>�h�l�Q��q�( 2��/F�ٚ�CO�^=e}��#���%�<�.�~ p��Ǉ�g�a?�яlذ�ҩ�\m��Qܹ���kW�;�vx��4 �L�dA���#(�y�r!yIՋ�
���ۉ'���6l��� �xU�a0dDo�Hɠ�}��G��}��s/S��n����SO���N:�D;��#l�����F�3R`f���"��=�k��؟cGu�x��ˮ;{zY��a��z�z�b��>}zI�ݥ��IJ��e�r�ќ�_?��z5�j`��; ������+l��i^�# �^:�Xac�Ye�~��}M��9g�cg�18��Ͻ�A	vy�l�1#ya-����4��? �et�I?�b�Ø��ʴE�;������c�"�)35�l:Tc������w�� �]';u�S�T˨VAQ8��v�6h��N6.���"��5Y��ɾ���y�t���lO���T:~|wG�b�G��N*+td �Y#[���۷ .]H�=א��$7�݆v40�%�N�O>o��jHk��իNF@��*W��.(��S�Ie��z�������B���"*�X���ch�H"zL���wE1��א�_�|*S*����J������姎C	�Y�e�Q�y��^��ZNv�W�̴�`%���z�U�����z_�Q%C��`8��k9xV$<`�6��e
�<��X*��.�jz%ov5��
��OcH�p��#��&����%�_(�K���F�;�F` �4F��ðU7�\p�a�<�զLM��TF�ޕ�h.]Yay�C'��>�.����}�\��tB��B��se���(�{xN$��L˶�Z�M ���gg$.�(��˗)E1_�܃����1Y0�0�G*?�����X8�|	kM^�D�L#�|�k����������Ce�ց����e��s����^o�M�<Ձ=��A���Xg*L}���}�K4%7�hJ���^�_�xAZ�yEVU�h��l�g v�J�_��X�Q�w+VJ����@�⬪��EK����m����T�4[�j��/���ل/&�M�q���}`o������Y3l�_��Ͻ��=-y=����/����==��}z�WS�ٜym��L+��K�Hݳ����T!�4�� nLĨ��\���!�H#u� Z!Ý�Gt��U���iS������W]a'�|��@����C;Ԏ?�8����}$��.K$�Ν�Z��|����F��]�J�ӂ�Zu�ʕ��+Sz��`�ҵ��2j��4���O�K?�c�
��1������{o��7ۅ\ࣤND�z@�a�L���m��ɟ�W�6A�`!�_��<���쮻�	Ʃn��)S'��q�=���O:ar�W����l��Ş7�﹗����ݔ��lҤ/m��肅����>�_��=��?��W^������o_{Ħ
|��M��O�[��su�&��J��,�z��;���]oɆ�Wؖ[nn7�t�v�O쑇��8]�������������'}9Y:�2�.O�����]�8�N=�,����'��9�f��9F��	��{�?l��֭kW�����>��P�𹟡�Y_��Uז[y�R�\��w���
�ۢq=g:5ד�0a;(/7ˎ?�;�'�ېaCl�7����)� ��
�sٵ�p�L�(��\���c��.�]�v�>0%��:wɷ�Namf��7;s��P^?�ϧ�����~�C�ؖ[n* =�:�t���6�l=��eKn6�<��cl�M6���{�(��C�����g�>q�����:9���A1bϕ69���?����&��v�Ω �e����}��(
=���'�lUD��bs��=Q�����e���͊ )R�M �wX��\�,��&�$�zq1�!�3�����<\
�q�K�MO5��ȁ¥� &�����0����`�-�yG�l&���n$��J+��h%�q� 
O���&SL�Ê��z�8��D�7Ěô6i�R�_��6D�4P.����7�E�Ey�"��9�{�$��c��xG�/PA��s�G R���Q�8z��kJ8T�i��-2k���w��{�Y�V�g�,2�)a;찣�GxȒ��ߑo��Z׀P�����G�C�R�6�"^�0��Nn�[����0����V@!<�3L <�f�#���1��W�mƌ�� {��9n����S���k=�&G_|t7���0b�&a[q:>��x��JZ���G]��h8e��EQ�8�C��3�B��!�����'#G���]�S�~��_����>�A��o߷��ͦ
/��� �+]��jj���Q���qUoK�.���]�JdH��^a���/��d
���[���_��1��}9i�}��g6n��6a�g�������Є���W_������;���+��u#w�q��p>҄:1B}��wJ�S�%U��m�T �-\&���p����#�O�����&���@��v���t·�|�.��2;笳�G�n~�=x��b�%���9OL�d֏~t��d�%�,G�#.2�>�NMQ�YdU�ַO?�����7@���ׇqT�^}��e��~�iʳ�N�抇
�N@m��
:����A/w�&�s �.�r��1ϔG� ����G-!�C~ȓ�d�g�N��
og(_�����T�;t��FK�̚5��4dp_���I���� �ܩ��QVX��h�_n����n���[�o��l��v��qc�h� 3 qٲ�^�`M'�33�)� ���������c�+���/��>��c�` ?o��&�.z�W��!����v�A�Sn��G�ſ��]p��v�����Kp�
P�~�z�ے3�3�>:��ԙEEE�t���w� �e��%C��R�A#��
@������*�x��쇢h��FH4�R�F(6L�A��aJ���4����8m���ٳ��� �>�J��3�b���3��p�|�� �H�#���1M�y��H	�����{���x[��51�*ʊ����i����ީ�oYa�<�Mx��#���h`����]��#���ߑ��=�,F[�C9��#�H����o�������D�9yw2d�w�^0�0*H��);���=�c`�;�ɰ�C���������Kd�})�`��dX�֢����Oߖ��ӣ42UЍq�y��Ǵi�\�態5��/���~p蛗�d�i�����/���F<�~ �Hu��o�F�g��1����:�<��b~&�E'�rI�3,O���(��/��~v�qv��Ϸ�������������ӎ;���:�J:w��$ u������?�֋.��~�ˋ�SN����x���h���ګ�l���7�����?(�9P~���� =;��3J�;HϹr衾�ȥ�^jMM6x�`O�UW]�8/�믿��Sd�eآG dF�!F�b�����ʱ.%�m��Q�Y���_/K�'�yQ��s�9Oi���p�	v��� ���S'�ק��`0��b���&|!�7�ʈ�@',�W���ga8�tS�~a?��O��Cd?���s��v�]{�5���oW^y���W����Ǝug�u�-_^��ZO<�$��"��k�'�~�k>�W
��[�	 8��8�l{H���+.W���b�%[`���{��ٖ[l�S%!��[������B �|�|E�𻭲M�ᏺ�)���z���ڞ���a�d��&��F����Vh���<e�����<v;���v�e�o�ݥ��?>��_o}�K��ޢ�.�T`�x��[n���B�dgw> ��o?���@�tt��6�C$�A�{8Lǽ���}T}����?>g-�uF�r�Pf�e�Q)�e4�� ��i��-�uLtb�A#�eBubK��Nk=����R�� ��i�P��F9�"m�B��2���V�� �^���	�р�xq��~R+ �ј����6ҥ�x��-=W��2�kEiih0�<���j�����ZF�b�FqMO�<�r�c��,�+��A��R�3珫� @D��!\a�N 7-�"o���P��S���K�w��?%��OdI<��0�@|���s�C~E��F:�|b�o�FE����"�ٲ���ΙcSe�(�a��/�@��!�ƕ�048��uG�
���)d�t��ݻ�zz%�*��+����>��]�������"}*qY�/2`�d6f \�3-����N�7��O�r��λ\����Ô.:

�$�d��Ƭ5��aD��� �{��'D>B��H�W�% V�u�(�s���8W�H~����	���X+�A�Iy7p�@1b�O�Y0�O����ns�ۡ��>�l�ا2 �}�}{�����X�����;�7^��{�}�������56?���^��>�#�h0������Ϝ9Gq.��ˬT��˗���lA�Զ!����v�mm��Q4]|C
��a�e5n��"�V�2�}�2��GLj�Z�)C����P<h���;P�g���=@�����q�����͓N<�N;���-���n�ï ��.��N=�T}�ﾻ�g:H@��Cs��{�ٞ~9���̙�}��[o�k���������~e�w�]�����/�.��~s���������uF��LF(/�	L� �u��v۝e�K?CѕX�(��-��!���6v��{����5��O��x��.ޑ�����y��r�!#dq�:n��P���	���y8DW֡=��c6�ϓ��F�MT��e�b�M�>�G�V,]�mH �-Sz݅g�0a9v(�5g�M���|���4���U_]�u�>�N3�4R�55�y�O<G+���^����I��a��ѥ�z��e���Vz���'@����}/���^S��RO44$2b��N��j��Z@^xQ����7S������1OÁ)-Ѹ�b!��s����(��ʒ�^a��J$~��#��E�>4�)�O��o�gz�ݦ����mP��ל"�ā0t��*�0��z�p��>�CE;e�7�b�h���Ɛߌ����t���l�Q��� k��n;�x�Ml��v���č=����q���d�[��l��v��W�����;��z�!�%��aࣥW��R	��Ǟ�Ɓ�Uv���(Ώ(�ΰC'�o��^/û{�nvЁ[��j���>�A���|�)�aX�Cz����g{a�=�#m�����>n+|T)�o���R�M�T�~�|����kj�}��-���w��٣��A�*6�ܓ�L�;ڣgO*����YX�nLL;">��+m,��XF|ܪ��n]�v�)PĉAD��8�I�G'�{��w��r^Ա�r �vi\�gP��è�_�Aq��S/=�
�s��-��|�)�Q����"h�רu����#�|<�^~�U�X/^�4!��8���w�Sx��+~�s��Y+��%�VY��~d& �a�OO�C��0�z:(����o�q��.���3x�<2C��2zG�Y��``M�G|�~:��`�A�i\����i��t��ZF�
%���B?�]/+/�i]����>-��Y\�V��>� �i%������=�؀�����wϞ=&���̦��0��l�UyS\,�S̶�<WX�Ú�y��6��G8L+#�ԇ��7$����(�Wp8o/;䐃=^��}�1����[��2����]�t�=��?��L�s�J��IB=�|8��[�����(�;�k/��������>/��{�ͷ|}�R_�U�#�sF=�\�兼0`�o`�c�\ɵo��V��t����ė�Q�C��<��G��Jc?�Ul��T�\��]�~t��n�~���ㄲ�T3�����םU?�r��.7'�%�����d����2ˮ���K�/��Ç�H�͜3�`G����ƍwp���_q�9����B��W�'y�ΒL���-�EK�/�i3�x�g�>�w�����ڝW}�4�=��/����<i�=�����K��+��^z��}�9�.7Ym&�22F�|a��[z"�&��ڲ��񩅯���e�p� S������>�z��W�]�R�G�Z��ڢ��7����8[��R�gȒ��G�C�C��D��-)�ٚx���q�NQ���䯶p�&�l��k���0�y;����hN;}gT^VQ"c������[o�K�C%�]Q�Q� ��F��hhpO�sO�J�=9��b@��0�k]�!��>�w:E���̣���6��i����o"�3�b�i��qd�!?ҏ��,��ֵ���fdj�s�<m;�����o�-d�2'F�66���ʰJU~���N?ݧr�(��k���^��3VPT�</[���$A88��U�\��'c�f��o~�[�����P��)�[z�� �V�g���4I�7�x�m��vԑG�[o�&c����>��8�+��O��nt�'j�|�r��z�Ѓ�؀~�|����|B�C����5�h�A#��$�^���a��<U���y�X�j�T�k�=m֬9ַo?���]�hW*�?K��H�I'qV��W�]`g�u�?�,�䛦_�;�YG 8�tT~�E��.X����lζ�W�4���#3d(�g��^�+����b� E�"�.�JF�{�a�K�X Ϻt �t�N\�1<��O>���)<C�/i2ԓ�]k"<dD9; V���m��z��|����.#�n��ܼ$@�)m���,�~!n���u�Ң�*�8��Kz�7���G��I~���f�`�I�c9�������)���/v��/���S�֘�{�zB� �)0r�e�فd�<�]�w,�GGBS�7��a{��~�%�����������K��(����F���qP��N@*uN��]�G��ւ�F]F�0��+�b��]Ǣ<!x`T������Lʺ��vʁ�%����3BB��m������!�<�w���~��#l��)v���ٟ�t�������_�1G/C�m�?��]����:�|����Ґ/�
�az���\�/:��upπt@mc�c'l��VW����s�͍��b���S?5��<�8������2(����z�LF}��ö�Y ���C�:즛nT>��%��%�G] ��CG]XVQf{������;���H�~��Yv���K/��g`�+@�|�n����D�a '�t}&]ee+�~�^�{܅Í7�p�ΰ��z�>��C�f�y�2�2�VU����|(,��2���̠��N�VB����vmQ�g=F+*W����Œ5v������
?G��	#�aT?U�#�<����櫗��f =��K��3LO���{��;�Ru��ן�p�\t���Q�im��Fs��;���<����vS����zG�>�)\����RAPR�p�K8��� �jh9;%�+�lc�U�z��h8Q�	2��Gj�Y*��+G���M�ߵ��kԒ�5����PR#�KH�K���i,�;O�:Yht������ޠ�ɀ��(C���1�@�gӰ-qYy�/8�1m������������-oy?v��>݂m��{�=���i���ˈ�1�0��'=�|���6x��O�ћ�����rp�&y� a$��n=���b%��=��}5y��/�����HG>�=�wб*�$�lT��iyY��8p�Ǡ�m�>F��*:�.I���Q�S���eUU�������x�~�_�h�
����ry��O�c��-��Ĝ��xf�?�
�	�07�d��2L�'����g�	§�pz��m���>r	_���YO�*�l��� !���[��Z�h��c��<��O����l���o���/��%�: y����A����q���i�fJ�	=��~1r���鿑-:�~;��9�� �/�z��;0
3l�a_�Ϩ';W1ݱ��R��9��Qf=���� �q~�w�uֱCG�b�-}�y��s���3<Nt�G�7�Xq7�(�l��e}UV&�`ĲB��[a���:�����=���ܐ�,��Y ��a�2�D�C(���.n�4���I	f4qE�J�2u��.���'�& �]�v�^={��A�td�-ia{r�Nf4���
�:$� �:�y��~����d�4?�*[Yj#G���rsx�)~ʕ���5O�(���O�����1��Y�%饮U]�����F�z���8��Qɣ����[n؉�2W^Q.�@��#�r�Zu5�/�z��ձc����3�vv�1X�'>ت��1����"�1n�@�@Yb+�����ж�zK�'~��g�u0��L������ŗ_�2K�r����k�6�`T�5;LYct�ic���v�t�9�t�ѪXnbY
��-�� � �XF~�C�xX�Buݲ�}�8�ƌ��u�����
���.]�	��+}(q;�w��9����xp�T��c�/EP�$��O���
��1���c������v��x{���������mxB�\S�;�K�^Ǩ�h���J�^L%�5;���1��6Hu$e_|.P���K/��Wl��������һ�7H�o�@���W_�b�m75z�#HP��"��BIe��?L뉍+�^�u�0~���8f��C���?*�P�x1O�^�$�b�9Oz/S&������SE�zZ����O*����T8�9�`i���v�-�x/'����sֱS�9�9�|K�ܑ#��C��K'7N_~�E��d'�x��q�Y6o����~g�~�Eˑ!�ko��$-��+���N?��G���]���]o� ����[�\�I�B�F8��H�gjhљi�[����W�v��|T��W^�a��PǆGm�W�a�#.Lhh������=�}�<`����G�O>�ST���0���c��G�ﰃtm��������]v��&� �{Ͻ�6���&�y�J1#���ò�R���'�yf$�!<��A8�%���66�%�%��w4�l�8$�> �Q�##�ځi��;��� �����=�65LC�C�=���ӓO�h^rz#<����!����a�ʰ�|4��_�WZي�	^�]���Muv��{ّG���l��Ɓ��@s�#'=�LEd�"<qX,��/��zԢ{a��>��
�i;�(��?��E҇nF�����45u���F��H�;�><���u|ߒ�0�#Yad/]ʁ�Mӛz]Jlh�V2��s�=׶�v{��2��/�8	�2���Xgw���2�Gv��cX�@�ӆr�LM'q`�b����idW_s�}�x l�CG2%. `�����N   �9㯃Rv�F��S� gD�8 �7k�HKHG�O)�&�B���K����c�ϵ�_��N7�UcJg�m�r�'繅�`С����|�|v���A	�G#�N>�iTc���z�/좋.v�ĔYҐ��r���j�c�S~w���+wˬt��3u���S��	,1�����#��	�J�)���U���z�q?�霳ϵ[�v��
t�2Ǯ� t�˿X�s�|s��0Ŕ:���&��i���#v��������{���T�y�e��NxڛR�U��`4&����Q�=��[�&�ll�=%^:���I�O�.��N�N�FcG�p>R(o�S�i�3¨#��w�+#ɣt�i���(�42�����';���ܛM��K���?��ݺK�"(�p�n��=�qQ�y�r8���N��B��f�g�8��^�`P�d�|v�����_�j|���vj����ӓO<5Z��w���O>��z�u�06FK�
/Y0����U�lyz����x������M7ޠ�tS?}}�7�K/��q*y���*��-�J�b|��G�_F͗���&��&�� (\��T�qANrz�YUQfq����B���@Ow�m��e���0&��!�&��{c���?�{��{��?�@����`�5	����+/���$[b1B��|!�&��S�.v+ď���+.���:Ӯ��:��%����:��-//sޣqL:�nQB �s�>+#s����?�Y`��O�=���N����&,� k@���"'=�N`���s��W��u�e>�2"L�{�q#�x�E�b�ײ�U�c�Ǭ�8���m��7�?��&��׿&h{�쐃�)Ӧ�;���ݧ�3 S �n��Z�5P��T�H��CV�*0�
eD�)`x��#��s�@D�N�g�#6�z��7�يW	��c3*٨t��A�|��+n������Kz�q(/H��2��9T�\a���w>.���J��]��|ZY2m�2d��R|�~E����r�k�=���N���
[�~%[�G�"� k�1��E1���}_+����M�%���β��L �ȫ�K R�S�hÍ|z����ǠDF���j+z��������e��cE�r(����"���8|0zؽ��}�9�o� ;��|]PMu�����y��npX.���OZ�ҥKl���^���q�A2ċ=oWG�~�9��M7�dÇ��N���P ϸq���A춿�棣�'Q��aO>���p�	J�b�w�}���+C:�N�}����;����L32UU�ۂ�}���<��|`^��������j�SO9��z��6t�(��deYi�5tRmH��u�u�t���4 �Ǐu�?�@����AÕ�h����|��$; 8��Aa.�{���"�;�z��6�T��7��6�hc��?{��Q@q�1H�J4V8#,���  A���t���C�e�M;:�(�DUe�]s�v҉'�<)3gͶ#�<�>��#����Ų���D� �����b���3�s(�
?tx��3r�#���Oz�Q�������}7c�����Gѣ��|/U^�&~1ѷ�� ��|��� w����T唓eL%�>c���,��SfΚi���=����y�u=�Y>��ӏ?P���Tdn<�A�A[�s*�Xy9_2B�k�q�fA��8ũѥ������شzҖ�� ��TQ2B�U͔��Y�o�}���g��=���C��ĉl��in(1
�t���}j����j�g�F��ֽ��ȶ��
��_�3�{�"�u^H�;�%�%�)��j���i;��I�Ԧj>������	��г?l���vc��S(a~���Z���s����c�, �<��?������B�Qww�Sw�S9���Sww��R�
�*��5!		$X����}����p�=B����y�}VfwgggVf[4o峂���"Qf�A����P�0y�
�^�	?��c��C��b7a�e�!�L+�<A�2U�M�8��4��Î�u읷�ݽo_���y���YȽ��۶���/��n^n��բ.��i-�� ���8B�C�!\n���YY5��no�3�Y�"� \W�d?=�b��"hg����d���U$=��H��z�%���eH�^خ�4�)֐b�
.mM�!eH��"����Ch�
Q(Ox_�F��j�fQi�,��'�yQ^�OW�jg�W5�}�j���I���d�X���rT��:u�A���g��:�F���~�At:B����]���j�^L�<�M��J͹.,F�cu��@C߈P�ʰ���R���}�fʹ{��gu�凳oR,U��ʶ��]�Q�ޯ����o��I�tчᩓ&M��>٦N��n޼�
�E��6c�t�6�������fy��J�	+K���U�J��ƪ�J�"�*U�O��mU	�iVW|�Q�־C[kب�5��׊���5�N�4�G?Q�b��uD��l���6s�)oּE3;��S|��!�J�&�����~������L��7�~�����![�z��%ŏ&������%A�n~>J���ʡ��s���~��K�].�Z��~���:��m0E������� !n����B{���|��	�+���2��*u����CW��`LB�AQ��`�y�z���DzI~ү���K�c[���#�(���3##�bd��-ml�U��,/?W}w��m��)o�a�+T��g��2JH�1���?(0L��o�ck�2� p��=����kL�39�6N�3Y��������q��$� �C8�����G�2�����)HP����gx
��q�Ƌw����-[��$P9%l��8���ɓ�oܸ��h�4h��u�(ʷ�%3��0 �a6�xq�mӽ��u��b���;���!����~v��~�;��o�NM��<�m�(��"SH�aJ��xF�"�Z�ܪ�y���bڒ7
qKRt~ ^�Lɒ�ֲUk{���|��駟a�~2�6nb:t�s���8�:� ǲ?�Nh�ɓ&���.[w󕟆��5�\m�?�طy0����#
��V��R�I^��~���`����sAӰ�4�@��(pű��'��"	uu�ֵG{�vڱ�]|�E����$�����WX�������S�z�\[�ˢ�+�	����I3�wp�~U'�VKR�!��{�UO���xq�=��v�9����|	�ͬ<!�G�؎���ᠫ�> �q�mT��/_�[���6B�5R?��D������G`!=�/@"�����'��V��[�[a ��C~��O�˞R%��By�@as���𯘎��� Ly<���8S�U;>��@~S6�q�S�6��t���mh� ���f�]ʬ�hV�Xw�i3�c��"�A���Q��w�3���������L��2!�P�gV��r�j7ӕ��-�2pN�Uff��G��vZ��0�A/��s�ڶ󭰜��*�6]�23�l�7V����f�6q~鮻�GyR8,�?�a�Z���+�Iٛh�q��z�mֶm[�'������oS~kկ��^��C{'hEHA���s?���_��ټys{���O��d&�Z�ha�쳏�	������P�m�k���.33�0���-X5d�W�e�(�*"��w,������p�+e��|��Ζ����>�,k߾��X�>�R��X��6�C���Q|�p���hw��6F�!_&�8O��#�+�>�Bx��	z,��'C�����+�>#>���J�1AD��n�%[����a���Ï8�}*�)�dڄz��pn���)�e�|�����gg�q�UE�R�	�&�]GÇU%#/8&/���!}p�=��p��y�~P�����1��'Ce�bz��*=Px~#���,]Z���ϓ�� �y`㔲��Я_��O�~GӦM��v���Ob�sS���� :gt��W@�B��ﰣ=��c���>�����{}�\�v�}�0�SO>�0���D�Ei�?��߸�c�1�p�HN�O+H��b�ti��m��/����)��b��z�� u���3�Cf�`pG�g�d[[a~���}��Ǭ}�N�׿^�)H�i�r��
�`)�q��y��
�M7^��6�n����8Q�q���(l���W�$�#t<���R�v��t�:	�2���8��35I�X+���M���nU����b�~�

B*ep�Q�����ꉁ�0Xb*^Rh�>��]�2Ε`u��h ���0�A��S�+�M��,�O ���2�	�:��JE�v��F��}K�@[x��G|{��C�7@���ܢ��%�K8�<	��[*�ݘ��U�IN��L��]?�u�Q	�3`|`Yi�����UP
Qf��+���ؾ���a�w�0r~�ZU�n�ٖX=i�o�cuC�;�g�~��0&ؖ�����E4B���Befe��(Q�z�#"�A&��\Z���`܁�u�W�"P>ڷe�Vv衇��A_�2e��ù�N�hs�'��I�H�����_h�3�}��9s��x2�o�������w#l�b�!B�>�h�����]�`�u�$�F��bN�����Q �i��Ҙ5s�����/��E?��83䕝�M����1�Vα��H
�J(FnC]�_��8�(}��W����R�0n�
8�o(��#V�8�D[G|��N��.�}#2�/ېi���MJx� O���ZV;�UM�f�[B��*U�3���l^I��T� �D9('��sQ�"�5$��hN% >����i�}�|���1�p(�(`�ٙNCL�qwwXq���J	���ԩ�<&(0v��M:�p��7���x�o+H|�)�ŋGJA:���nߢ �I�?�C��&��EEE����g;���Թ�%�3���Wt�6�%K�y������O?��c(Y�Tt����z����0�dAt*�K�ɻ2���2tn4�mT�o2��311w���!0�[�j�(��JԸI�g�s2c�u�?��{���K!�z,�`�j���ʯ|%b=#�Z�($��>֫W/1b�}�՗b��\��m�Li\�3��0q���e������s/kٲ�[X�4q�p3�-�"�&���"���V����_m�67m�d��S�WO� H=�U��e�ώƀ���AUw�mXU<����WϞn����^�-�lmC��JϦ@�!�7����q��l����7[B��FYVT�M��!h��C<���QQ����BEB��|�p�yz��	a����
mH��o�JA�Oe���'(�a��.<�A��3�5��Ί'���)�%�Ap�o�2��{�Y�*������{V�Z�n�yC߄��i0Z��gب�̬�u�!y:����7w�Ō��Q�񸣇� <���(����AہKڱ�����z�	��Of��R��Y�@��� ����a�C�/�'�VM�%�:��ۡn ����R�zo���*skgÆ~gcǌ�v�ѕ-�r��������Ç�����cF��qc�٨Q���?�b?����U�����N�����[}��G���/L2�D�C�F�����߰AC�p���la��u���L�3��?���7�m�7���7��KMO�Pb�����3���5ځx(T�}�&���v�=��	o�a�' ��ޖ���ą~��ڢ�Eae8���r-�6� G��4ԩ�V�S���`x��%tQ9�8�� � x�#}�'t�x�;�	@�Y-d�c"�>�+��P������Pv�7N&t�A�{��3ϰ#�<�?�p�Q:u�~�!�i�s�ݺmmGq�o�?���ܰ	�Z��-�������sĳ"��
�/��"H��;ہ�7�C��[o�m��?�'{��(���?^�&�dI1�J'��0�dDG�Q D�̢�g�ycB@�neK���<����H��!M ��+2��@Xgΐ*w匣<�T�n(S����O�^��`�x�b0�E��� ����r�A�|�������u�S�@�ij�%�P�.�Ϡ��/q����α�v'-ʅ	j�0�0����P��[��)?o����2�38������B[����K(w�v���!�T����{�xF<H'�<p���'L���0�3O�!�\�i/�ʅ��v"}�e���8S�#>ɏ��N.�q��?��i��(u��cɐ�-9O/����*z�+]�\m-��IA)(!��g���ßd�/��Xn?�.�d���K/�-� u�<@��m�Nt�q]�tq���5�Ȥ�M7�d={��ҵJ�J0-�KR�\(�cT8��B�xʱ*@��>�.�%+�
4B����.?���5=�V�>q��Q��>c�\�<ڶko|�o��N��]��e�������-� ����/�Eu	[Gq��q֙���ǟ9�Ԯ�m�]�7��o���A��w�}-U|���Ř�[�:u�lmڴ�Vʟ'F:�� �+���vm�[�N���c,cv�{g	����je�Nh�`r%)����L�ʬ�+M9R�rj���N��J���-������p�����������R��I]1��
z�������U�&��q�.�rq.f�6l�24O<���)��7l�H���:w�b��N<;v��u���f�Z(�F֨qc�\�%%�]ݶ�����]���c?�ط�W��?�G�����I�=���~d ���||x�O������8w��Ίu����M���cb:ɀ_��\�@�\�p��7��Gi]:w�V-��kټ���L�:G	C�ؾ��7�6�Zz�޽z�q}��>ҪU+�3��z�������?��/����Zcw`�[�O�כ��	4��@�BLj��`e���;;�  [�r��ط0�+*.v��Q��"ha�2��cI���(67�~p��D=G�#Í�Jԓ�e�!�t �~1(x�M�3�żb �0�B��g�4�S> ��l��5�Ҟ�+�j%������o��<+���ii�"  ��[4(?�A_��0J�3�E�o� ֕;����V�.��{����淧A�<HNBo|��Px���#���,rǻ'��v���o��~'�M�����}�w9hM�`E��h��:qy�.~��;&��,���ַ�H\�I?e�h˖-�o߾֩�Vn�a��e��P��8�t�e�]<C�`V���[
���x����jat_��9�'<�L��s&��A��wXE�ۋ����^f]��n_9)S�R.�/���� �@#T�%�-�o��Px`����U�[n��~v�$�t�	�=��c���Q��L��h���R<Y�AHE1A���t����>"�S����̘�CIyX�\-����-��[RB�h��X��J�r/��j��5Τ�
��B���Ψ����#/�
|ň�'�UO\�*��Go�`H \�.�[�Ly/��ĥ=C{1Ŗ�
W�t¶e~s�RP�0,�L|�'��6<��)�ԩSm欙N#q2��G�"��?�Pb&��p�#���Jy��c��㻧�HcS�p���xF:�(J�F!��F�is���	�ȃ�!ߊ�H�J�ۈ3x-�7��/EV���y*L�H#����"�j��0��āe@y��]�.�Sю��[U�o��LyUR�-����z��FAgu�T1�ja@(K�_���LH������f��>ls���QE��Q��tar��5,0~����O���l/��
Z�����gp�� �0�C�@r�ry��f��jpe0!}�F9�7��8��3d��0�,\TD�!��X�~鳄������@����#Dz�I�;}���s��Z�;:��(•:x��O>�^L3�';��ݿBy���_����
����K�cЅӬ��
)+�� $�pN��Pb�ZUː �ц7�|�0\�"u��[�^��F��B�,�B	�RݕY�7��v=|6T���������PZ�YY[�s�~$��(o��_!A����~�Fڵ�z��-��B��4`� ���+��+��G}ƞ{�e���1}�[
(b���R��!R�p pQ�=(�$/�zY�cR˒�qg�BlCڎ�qRk�k쨦�&�23�\e֔_Z�[��˩^���zǤ4��ki#&�B�i��D~�nb���i��vQ����^PRp����_Y��)M(�˥���ry��e�o�\yB�^-���|[\$E�t��W�W$�(�O���d�hڴinr<�j W|�z_�T�Q��I8��c�X�d�Ɵ��DGX\̇x<7�7�2��I�<�9p�E��r�t��D%��ˏ��O�\���w����B疴�ejPf�&]haƬ96O�y��\�6c��6z�=��K���|U���ĩ�.���?���O��w9ʨ�P�ę�@�[�O��[`s������P���85l�t8� g�	�g֐����oֵ�6>�
��v�Ņ�
�ڙy��}&�3,��[��_^�>���o���'ׯ�;<��&a[�!�=*� �� 2�8�^,��������w�"����.+8���3a�`�:��x1=��6m����L�/�Q^V��
y���A�ȷxI���($�S/~0[�
�e	4@����d��*�_����-�"�B^6��8���ĉ��l��5eN���9�a� 뜜�!�-���ڶooݶ�֭�!�r�M�{>��ֆ�~ہ�:��N՗��J[�W�)H��Z��4L,�6��w�S�sa��/��Y|��˷�~o_}���	"�}��׶�fk�C	)I#	��۶u>z �����clT �)k\1����$L�G!\ ���i��L�1����@Х��r�ʫ���ږ�UG�F��+���yp��L�*�#��B����r���'�W���2�8�q2��(I�Ǚ#x3�iiR�OH
�~÷��8���I�J��I��@���xR�a�1*�`J����ۤy:�ЖL��YYǡ���}y�'�͍󭁆�2M�u��v�:���pKi��Ħ@lS
D��� �8��"�jڨQ���Q�9D~����bY�������k���.����{���-��j��w���#<��IYB�|���줓N�SN9�N>�T;�ē�뮳���{�cP�۫�'��Q��2�g ����F��TP�ȱ���>Uu���[��!�0����S#-Uj�=�ܳ΄��g_g>X����^��s�QT#�cp�o�HOϲ�;�N>�T�$�L^
��_��FG��8T�)����Jv�3����g�[���P!!��%����gqb�O�����0x�p��V�4r���Ua��C��&��̕ ����z.�×��g/��C:�;t��V�0�`N|��¾�Bp�ABH7� l�A?:��'��^I7==ͅVM �(,a��A Z���bx�g���Bݑc2�Ut�=�y�
a�y���w�۷��;4S��+�Ji�+�ܑT�?�uش�f}G�����?�q+˫bQBXx���Ejk.J�;���0֕l�V��ZJ�R+.ZdK�pk��5���c-Z����ٳg��ɳ�>��%p�	Z��t�0��=��Q �̕����s�7p�v	[�E�ꟸ��9�_Uο)M���~��b2}��0��@��_��I�^ۻp��/��?a�J9lղ���y֢Y3_��^����"̇-V"���l�&^G� �TW��j� ��j��U���u�����"!&ʧϜj�α�e+�� �D��|)KS]a­�YeӦOʗ�P�w-�Q�͞3Mm8C<b����F�sԏ7]R%����]^�u��Gl�M�7����Po3gN����ۜ93U�|��3M��cd!W���:7�!0}�|�2k�PJf��~�|�	���G�iek���d��Ht�5L���������U+,�0�J��*��6j�8��l�c{b��Ha�z>,�eS&��1c�X��B��������rUU�q�B��k��V���q�!�'��s �ĳ�Ŷ��8G��?c{G�MYQ� VQ�P��JX�����7ڗq�o���n�U��Mv���ڽw�m�G|�z@q��c d����!C�}�ر��Ge�0�c
����|�>�N�:H���-���$�s�sm��5$X��\�V͜�̌�1�5l��;�;ap���W3b�:���b��u�9R�^q�Y͏����Z��~�
_˦O�e?����j֦uKՀ�P:0�ƃ���g�`Bt��U�0I�h 2�ȗ�i$W�û�C�U��ʅ̝r&�M����d].���B��Lt�\ئ�R�e��0 �,]���/�p��K8���lG���ٵ�.*B����`X浏�ኈ~��v��s�<;;Ǹ�L���e��1�1��:g�G���T�U� ��ٷ���z����Jy���	͚5��4��U���`� !�jY�d�4��=�S
%�RܛMm��dWȻ���0���\��AX�u�4�pԽo��3��p�Y�$G� ��`�M����S^��7��ܥTQ['.[��6����=H��R~��$)m����bV���{O��oWَ;���9ٶϾ{�g�m��*���+��/�>��ئ�GmGy��B����J
gb����L7t�Z哠Z&=�7Q��'���L�A��r%�c:��קh>!';�c�<=�[ŦO�"���HɨQC
Gz��r��/�8l3:��ܢ�7�`���x�߭K��V�V�5�_�ڷkcݺ�գ���v��	ǟh��r��u�6{��u5^��@�ǹSF�Z#Z�ݶ
�п�+��X\η�9~�V(����s��Vv�}wۛo�n���co���=���֣gO+\�k��4�g�y�^z�9۾�66m�o6u�8˕R��^��9�ku�K9���d5�)��v�0e�Pʛ~��fU�����`<����ӥ2`��X
H��w��Kj*[ĖXa�?'��H�/�UU&���η�RK�+X\d%�K�I��n�h)+(j�+��v�^�Cb˨H�!�����S�0�*m.�^�r�UO�fݷ�֎<�(;팳�/���8@
�b	�����ܼy���l��w�����{o�a�����.��[u��w�]4^�&N�nc�L��7�rjgY�N[)\��B��?�M
W��	*X�<��	���j�)�G��U|%��Qvs���D�Q�?!~�x<��]c��s��Z7����lE��XZ�xIx���T��FBZ�i���Q�H��0��[��xwy)���������7c'u�|�J)�4�v���B[�_��n����b&k�`R`.��kV#�0�"�S��ԫļkJh�ɩ'�g�=�����+�����*�R�7��9U	�˗�ڧ���y���6��+����%%�,�6L(	8:5�8��Z�)�r.
X@dJ��<a��s�����Y��:�@*[	(�OYPxGA8c�-*�9�����P��F���3�b�lE��A�<��)�ps�3���� >��Ղm��U�8x�/ab����)=W�nQ
s��a�8 .liB8e&�#pbĴ+�(�B=E�� �d F� eJ��?��v��_��]��'!<t����y���L�6�v0�����;�`��׳��O��ER�.����z�^;��C�J�5֢Uc;��w��~2ۉ��~������Z�v�DZ�w�i�ϓ�`E �q(Xc��̚�3B&�'L���0���O��W_������c�j�i�/���,������"��)��*�'� �l�?"�3�?ݷ����.��+�P�ុ�f�ﻏ]p��>���n����#�8�n��6�֭��)�->q�7أ�>hg�}�O
-X0_y�mŕ�c�1L�s�>/D1����n����>x�Ϭ����N'������Ř�����7߰>}v�yR4f̘�vZ�1N��	��>m�4)H���*���>|���M�93�@�v�����xJJ�v��W�no���x������0~��\��]�����[�ً/>��d�����k�oك�g[u� e��m�ڞx�1{���v�%��Y.�,; �=�%��� 壈�T���V�y]�;�o�n&#P���L�A��Sv�Z��Bт�ic�,�<C�ǖ_-|ɏ�C�{���w<�XQ��z.����<����Q*r]"��3�����@Bc1�b� �W��1��~f	�Rx�˅�bB>C]�2ҳ5�6��_i#��`�%˭V��b�`K���o#U���믆H�)FXݷ0��l��U�Q͸�,^rV#��q(pl/�r���H�h���@��`�DF��+�O�~�$�D �Qgq���(,8�>�AR�irY+-��b��a��}��8� >l�`�B�8sx+J<�VBx��ξv�����d�BX�Y�E����w�h���^'^<gम����7�ؠA�Gh�Zغs �I�6��_�����7��S@^��'u�Mk��	b�Q���ꫯ�))�?,�~�M�1Ɇ���~���r������P[Z\dֶ�M�����Ǹ��7VK�P4��[y?�7Cl��6�ߔC�M;�ӷ��I�b�~�P���E�_��� ��>��s�vG����s��}���-��R�6�����3���T&+_ą�qn�;8�ye����V��tݪ�=�ģn6�W)��{����ݚ7ok��׳�q���F��Z�����+i����.
���7�n��E�rm�y�Ǟ{��p���Z�]zۮ}z��hg�q��w���m��b��νm�]{��?�w���}<W]y��b�{�X�v�0@��j\�E	\�m��ٖ��n�]w�]|�E֪ysK��UUXůW'ˮ��
��ָqS�QŚ4if�4���9V;���k��zo��z��n�Z6���kى'm\x�ee�h�ΰm�mc�۵�N8ƚ5i����8�r��7�&� ,�,�٢�x�U��K���2�{��v��ݻ�Di3�J�������-\�͑����O�q�e��g��I�m�h��L]����C1����N_�������7��
O�B��ַ?����uR�����%K�/^�8#�Л��]&�F��\	��hPY$�^$FS���8�#��3�a� ��g-���1�X.�^L������1���H�� _�.֠ή����qa�ɯ�x�$��\����X��ѷ�QƓȠ`h��"�@��&���A ƍ�Ae}fdQPx�41��PF8ډ�v歁.������8�:r��t��p25P��+pB�6�J�D��y�G�!�q�= N�̌c�a��.���3O�p�m��	n�hĈ~E���dE��F 	A�m�2�|���P-�i@�Ӯ�,��r��=w���C �R��0g�l����G���?�謴p�

�Ih����t�� �C�� �ￓ�b�� ����ߺ�>�~�i���8K�]JRX�;������~ۭ�a�����		&���v媠p5kմ����;(q�V%+BeuQME���w�$��J��Ο���ÍS�?��s�裎�s�=�~I�ǜ3c�SO=i�w�]��`�|��v]��kש��?l��J��U"�Lv�8�3�u�	�t����"֣�ֶ\c߄IS��?���y�mp���3�<]u���5�[w�h7�t�r�Q���;I1ឥ۾W/?���[]��X�(Ӷ� m�bY����v���Y��ȁi�ym鲥V�v��y�ɶϾ�I9YecF����(T�ss��Im�����-�i������r�q~Nʷ
���p]EwC;�q����ӓ",�&(�\��6���:]m��g:�[�9�'��3��Y�'��-�n-P�%��ӥX>���E�ܨ@;C��1��i�x�/����� ^�u��.[�O[����VU�0Y!&S�`+�HAa�U�^��կ+�Vb�����s<�1+A�>Xr�^V�,��-=#�#��Sײkf��́�<����?�Nj=[·`����Pq�<33��~�-�_��Xv��>�%2�d�惮���?e����@Oz8����w�a��3Ϥp��pV�R����d��LN�p�*O��lud��� ����[�[1��+>���:�I�@�4�6"B�c���b�,�/��&`]y�.^��}�c��pa��b�?mD�p����'y��	^�ȓ�!n���X)�ҍ�m�=�|�#G���V"��x(��3O~�o��q'|l�>�Gq#\|'��/���p�;�Ǹ�#\�;�Gxhቋ�p�+	'n�'��-�@rZo�	��-��./���x�hfQ^��=w�f��Q#C��d�⋯-/7`(D��5��J,h��r%�.e�O�hl?�&�!�+�p*/�{���^�%�ߣ�g���7�r�<�C8���N=���
O����e>����~���e�裏|�p�ֳ�q���|��'��@�6��;n����r�������z �)�VL��#.�=��N��Qw�
��� 7\0��������j��z�}��0{��Wl��!Xi�as��'�e�]�c�N�jnB��pc���"����aE��p�/��:|��U�m�=v�޽�󴧩>/��2;��S����_�G���h<-����z���]
�M7�h'�r�_� �R��N���H���خ/��q��о��ޠ4�k�Οg7�t��}�i���ߺ?�u���M�>�|�a+.Y��;�m��A�d��OlEY��2k e��K/�k���իW��Y�d����7}
�B��O�8 ����	[�Y�C�!��8��e�(3|��������kƣXg��b}�z���"��⸳����ڃ?jO<��]q�����_H��1�q�LH+��.e��=����6mi��B8�3�&��Z��@�[�O����,@�.E� �N��J��� ���{i��^|�9{�G��{����w��{��}��v�����������7����<����a�<��oqy��'��g�����>���㡇Ĩ�G}La���ۮ��:����ʫ������ޭ�۶kk�͓�D�S���\�c����u���mMPh�4��.�;L62���l�*��1�hvՙ��L���4��w,Y��803�bBݱZĻd���o�#uV��G�b�}M�J�����<�A�=����rD��a੾n���p�R���4@p�~x20P�:Vf�p��ܑ����u�<��y���˙@���\ ��˼~�+��Dp���a��żxO�������7މE}�֘T�EA?�%�Ц	��QI%ﴽ�;O	ڸhB;��;�x���Đa�ܯ���� �����?�EGz�H���I J<x�:ę�fM[*ϕ6l��ríx�R�M؂�|Y�͛���,����/~�d�>��g���~0x���Vb����#>��� �����=�����?���̠# �ݕ���z�NcYyR��V�to�(���$��ExZ�t�ǽ��]�g	s��?��~��o���xf�����Gy�y.i`����R�km�=����ނ�������v�x�i4�+���>�@\]�6mjg�}�Ƌ���W^�sS?��o)kݦ�]s��Vk|
�j���Z;�� ��kxI ���
H�} �X�@,'P�VMk߾��l�BB{�����ֲ���P84F��Z�m���{��Tᶮ��	���t.��%��DK����}�1�~�p��`M�ti��˥(c�=g���J��neݺm��\��Wv����n�E��.���J���G�L����-����i�Cp���r�ic���rT�:l��'�j6e�T?�r���?|�R�MH�����9/Q�a�*��R�e�x�(E�ꫮ�K.����?@�W�5n�D���� b����dW��� �1��r��������cl6@RGOY�6��+��Β"���֡cq��v�A���;oo}v����w�}G�ݻ���~[?̹m�.ֽGW�ҵ��l#שsG�ҥ��h�\L��rȶ�[�N�����X�&��>��>�<�@�w�}��v��;��������mW������SOw�0��LW.2��6/����+���m�*VERTK�)�%E���,�`��ǻ�	��ļ�����/�1uf�
�W[ �ʀ0>�%���`�@�3̌�\���R7+���`Ny8/�`W�F�efe��[�K�q��y���U�B>�i?�]��4[��EV��PuT�:*����  ��IDATB~k�,(\d����V�.�B�B[�p��b�u߮�_�	��A?����:�%/8G���u��*B��2?Ҫ,=��t*~�q�]���=�%C�M�1-�fW32YUIu���Y��G���.�!m�;�����Y�I�}�}��u�n�m�����
���Z�k۶m����m۶���ݩSg��@i�l�!MpbB��3��0G��<y�݋�LD!��3nפ(/F@&L�h�}���/ʷ��0�̱*�Rm��9��o��_m�n�����A۫��jGu�+/&N��x�rj[��ͽl�պmg^圛����9�KY���O}bpE�26������!�f;�˺�@ċ+��0-G)[�
tD:�OA��M�ӿ�/�#��ϰ�~�J���F�����k��n<P���V�9^VF�A٣G�6��<��ިt���� ����i�6$�J�@��,[u�l����ҋ/���m�u���ֲU�{�}m�D?WQ��_F�����&Dv��H���"�'�,��C���[�_q�}���I�Z��>2ě��� �@y��[n�^x^c�.�-Y�8oˊ~8��ܼ<�e�h��,JuD8�	D��i|��T���Z]�m�.]f?����i�֤QS�gE�q����αm���ww LR��fّGk;��ɤ�*�*VX���/�b-�@�T�1����.�;\�X�X�u�"Ee���S�N��#u(�&N����4-��3��6�aC�گ��bcF��m�leB�# �ٖ/�f��>k��XMf�����mʤI�H�	��b2Pc���ޕ��2��@o�\!�Bt�m6�(�oR�o�Apl�4�f3��l��'�ܮ�cP�sM�7u�@6����30��׫��>Ρ���.� � ��53LP���%���Tx����:�-�:��`M0(��4m��g�������N��O>�Ԏ���Ϫ  �l�.���[d�`�|Jf����1F��]2T�JՠQ(-ˤ�t��ͷ�P��_����Nf�Q@"c�kn0b�Y��-ZZ�m���ٺu �~��_��4ފR�""�y�d%�z>��s��_��o��3=�z�4��^��ڗ4����o��!�:v� T�.��<�~ؗ.H �a���Aɕ�ugG�q��`�d�R��V[���<��~�=�h0��㰂�;�oٔp�@�݂�	���w������c53k������2�h������&�}c���2��ʁ�O�U�� ��O_���X2��Vtĉ��-���%�u�2 �#<a��(@3��Y��E�P��,��B���Q��a�"\<��.�p<���@��,O���7�Kt��(�a~B� _x��	�<��{,oL���L=���-���VÕ�?nݭ�����|�8�/Ji�<K��/t�p��y9� ���� -�k�P������s�� Δ�2Q�q��Z��P�e���z��S�'CVr�cߣݸWg���~s��{�i�ﾻ����k�Vm�ʜ����>V>h��aѾ�A�z����ҜP{�����f8`O��g�~��[�ꮱ��e�	0-�BA��a����:+3ۅT���l�.(Xd�T���p�����mL��Xp@5��re���λ���v��'[��¨1윳ϕ�=���.;�����M�9�=�H��::���ԕ[��`d&E�{͚�h ��L8V�Pf�����8��!���i���40h�'֨A}[��'�xBJ�h;Z񎖢WC���]~�������h#̑39b�et +�e��|E%o�]z��v�7��fX��v��'��AZw��=��u��˕��O=��{�=kԸ�]w�5v���~��s/�d��6����sN�|�h�z����v����ǴԪ�����ڔ�c�C�v�?��R&(Y�d���P�;ŕ1�I:�@���}QQ��G�cԷoï.2��(��-蘭���R��'?��?�i��b�C>\6��:�Hg��̞�g-Z6q:���\��(�����&�{ �^��߆a6�خɰ�x|��3���
�ѩ���01�z����O?�K.�bl��6N)[�?
3f�l��_�^�Jվ�C� s�m�ȣ�t���?�h�����;��L�8���P�7:7%LF���(��a���Ơ�a���]O���#C��\
� �f˖��3ϴn]�:���N:ɕ/f���jeb�H0҄�%æ)H�/���8!��c� |�QAB ��
�!ܿ���~�$�lnq�0��q�B�Q 9Å ����E��[JA���0�1f�D)w۴)�,-#�'�J���2{�ŝ*[u���̳��Y�V�[ZC�o4�K����'m��ɓ-%XO<�OZ���.��`����6n��'�z`����NA��Cq����=z٣�=�BX�R�
��8�\Ct�@M}���l�L=Jg'���P�f��A~�Iv[8P��(3XR����c�'&[y�+4q�^e@:��`���t��u�őx�)���ӈ8V4�pl���޴A�W�h W��6�b�g�A8�/��~�c�0aU ��Y0��Zm�&\�R���7�+��A��IY	K9\�2��O[���]��� ��|cz�Β�&�x���&oo���f�/-��	��ee��(S������H��!m����i�A���+�!~XA�
(����u�S��]�pB�%>��!��74��M�L)���0���\�%p�0a^*%�ܳϱ]�������n��~�~�ڦ��Y'-hPi�7i3y��_���M�<ŅL� ���Y�:�ز�|Y8�4uP.�z��к��Q��?yR�����w�y�]��+<� ���o��پ��g]��S�̰�Æ��(����o��"� :��{�,���fΜ�0G���c����簐G��meU�m]P�C�Ϟ9ӎ���R<��R*��觟~��k.�����_��^z�Ԯ��_���?�'	/��R�C�Kxw�]v�喷(�u�³�C���h	p(���`�T�۷��r���5��Ι�c�_�.[u��^~ɶ�n;_�:���_�~���fg�s��~�m�V=�>��c�쒫��㎶[n�ު����kv�ŗ�}O^|��u��7M�}����L� ��������`_���x'�ߪg|Yi�O�����Z�[U��_1�o2)M(-=�m7ܣ~����Rn�<d,�j���D(ϴ�N[St�6��&d�sP��L������ì�6a�8��Vr��;)�B�V�_��5փ���vc@Zac�������W�Of@���O9�3.���-
ҟ��b��f �]qE��c�XPX؉ez֨�Fۘ1c5��j��WD���Z�p��j��Kp���r�K����kmI�214	m+$�./���Vq)�r�K<|��uh7|�I�jhM�6�΍�Ϊү�����c�ݭQ�`)i�o���?�� !AauY`�@|�@R��$��i�0�|a�w^㶱���ܻ�����|`�A�(saň|W���X�+���
��^�歹+$�I1*p��l�7o��7F�LOs2�С�DUW=&�&����^�)� @[sI�/���6����$���Ͼ�������#��رc&������}ai+.M)�`�SE��O�,����6�].�Ehe��O�|� v�����4�Oo��q��c��vک�@
�M(q��F���^}Օ�L�
^NNMϓ���Bm��0�N}�Ob�*�qqq �>���Å��O�AAa`a�T�볧G��!/�]��'���TB���XYê+V!���`��Sȃ��qP:���(�>V:ɀc4�<�kh�rDG�B�70!�'������E��� 7���0��[��E�t�e�6�V��B� \7*��� ����kH�Z�-�9�b��؆���A�U&+���B�"�?}��h�(\	O=�HW�Tw��ۅ8�7�i�:�=͸M�4Q�|�]��O��X���Q��N�;�@0�T�o^�`�ou�!�w���ƍ�_|!���LJ�/��k�Y~o]��͜�7��ط��0[�E��]�`�S���h#	���JQvꔲ��F%�6e+.��~��ù�(]�[b���X3�ѽ���^N��:m�M�6�)�-Zx[AcǍ��m�:�]@N�]���^�B����k���y��7��Ek��*+ǴD_E}�X���R��t���K�h�v����%������?��Z�h����X���7�|e}��"<���1����T�ֵ#?�z���it�Q~��`L�7��NBU|{���^�;&6X�̔�?g�|�m�qđ���T�|)�̝vG{�v�a�.&��j���Ǜ-[��?ڧa��6o�L���W�.[����������(��R��~�M���ެ��m�	�<L�09���U��:.�����e%�S�RX�"��M�ҩ�:�/e��5jTO4V�jf�?I��g���-r1�j.�sR[sN�2��I'o� ���s��7k�DJ?iղ�M���{�^S��Ͼ�1�vFI����X>|?(�qL�ܭ��*��/��O|��腺�L5�gϞ�i�-��ÿ�R����Ϝ����o���a����}f�@�@	�f����vm;i����DHp 0L����)iᇰL2��F�h����:>в�e��R;����G�=<�w����:K�w��Y��U�2O?�m�P������?�U I1x���4��T�U���q- a�f������I�oQ؃�1�[f�֫�a�h��ѬYK�4q��5�V���s�r�ldyy	�P�J��j�)R�`�X�"$�����K��Kn�k���7�a�����p��/Y��=�2&����5(r�zfy��
�YV�8ۆ���7�X�v���/t���AW���%�"~<p����(�.Z�X��/�i�%B��c���0�������"#ۊ��ZKZ�K��˂1�OL����rC�EϬ�����n}�}�v6x� +e�Ȭ�uq%���Ч����̋>�3�aU��؉G��WҢ<����=�u��C�4�<��aq(����"� b�[(w���6u�"M�^F>�S� ~ �by�qI�;u�o��yQ~~�|��0<�;�'yD?�ĸ��$��=R�l�ae��"G3��$��;�۴ik��7��z�m�B�{�'ՇX��
Xh ��	>�eBU����H��N<c�杺�&�"ά��S��� |'͠��jn�3ML� ܟ�?Ǻ�V�^8|϶�L_I�$d/���z�M�e�����X>Ls��uo�>m�uݺ�|=SߤC��uQp��C�o�[5���"5n�߯����D�|��W6{�,�G�G��V5��x�v�-���C]�n-���*�ow��E}0�'{퍷��ϐ��\|���Oz��U(	@)��p(F��ӱcU�f[��w�^R&ͷ�B�����K9 
��f���~��	'�dO?�����G�O>��{�1kӪ�� ~7t���G
�;��u5v�D;���U��^&D��CA�� h�luXQF�Z5E<7ӷxϟ7�/n�~���x��ǖ1vP�l���x'?�g�����P.ɇ6����u�*;˚6in�n��J�ũ�����WI���ο�f͚n�r�4� �0�k���#?�� ��`SҪ��*� � X��<��y�w�I'�4%�n��6N)[�?
S�M����~��o���T�;!��\BJ���ݲa�6i��Y͙#�q�u�'�C���qq���QKG=˗��7,�׮]K�l;��#=����>���<����&l��l�*�%�|���?���0(i�lm�@)�R50Dؠ\		\q"�N��'d�,f������8���~�,&��b��&+����5 I� }���z��� �B��R֫����ay�p^���5�G� X�cv��d�ծ[�ˎ`�,�V�B���/W���K�S��K�� ���KWB4p�2���K�3��c�9�Q���ǡ� 8�_<���-V�իc��~�u붵��}��7��/N�\���P� �WwE����FI� ���ҏ�%���'+��.p�}�'����O�q�S�c]��6�g��.D�e0�I�8|C�O�/����". ���#=�gt1��iIq���ю��/xS_��aI�w�"����b��D�I;*��?�<Y���pl�� �ܾ������/��';��#��P߾����g����'�)(ٱ��e��¤�1���M¹P⡌�3y�x��Ohw� ��+�"������_�m����7+���l��yv������`�9&N�b�s�:���V;�s��V0c~�'	��}��=0>�I<����v�K�k����ɓ���[wu��{쾛�r��R�����>��c{晧� �_�=����+�Y��Y�%���B*ZW�qq.83&�4@�O�3w���w�_��,��*B��|��{���ǔ��g��U�b)�l�,�>�[��C����Jڍ1��~ ��L���C)G^`%��:dE	�&�9m,�ϖ��J�(����{���.O�`�m������>�-&�����[l;�,Ք)S��EF;� ��W�ܒ�%���v�m�C�.]:��&�jTʹ�>��.���:u��Ԯi+W��衍?��Ċ�_��*�����.��N8a���'�-[�63������j�k�<�e!0��Y[35���{z9Mǆa����M
�L����dP���3O�c�F�F؃���1�9����]$8 ��0�>x���[8b�ɰCI�R�0��T�}S�X��?�Q?䬂�����չi�V]`5}�^#՟l��!��߼�J�%.�22��,"US|VD�k�=*��t u�#��`J��G�Hʓ�\�p<YU&�ׄ�Γ�)5U�TF��A���o�q7p���Xԏp M\�>����	�tQǔɝ�a��,Xu!l��:�](��S�К>�T.A�K���(���gE�����: ʅ�J�҂u�m���:u�l�ڷw�e�.]���7�w`���&����J��������l��W�Y3gHp�$A� ?x���;ٰaCm֬�
�F�`냫}�Q�֭$d�{���I?��ǲR~c@�w�KDw�a7R�J2u�@�4�weeu�6%^����x����7yb���Q�ĉ[�b<ꁴc���NL?�5���0�G��i�p�̸؞.&ڑ6�� �QY�tKX�8∋?y�? �H?�C}'��{taQP\I3��T���:�r�q��w��Ռ�?T���b)H��V6���h�4kp���fϞ��B����'�@c�`����ߜ�[�g�EŮ���%
��J�hE
a���(�hw}��|�ܫ���`�T�+�y�ѣG��ִ�m[�D�t����<���[o��L6���HO�클x�<@��G����ɓ'(�©�� ���g@�k\+�s\�-,,P��ҒR��
	����q�P��)Sl���ֱSGkݪ����X��;o��|���ҋ/�b�����|ŻU��^NV����3g�����L��+6�3���͚�/h�['��
�U��>TO��[�'M���Y)	+_�]l/����͎;���+������r����믽���9cxTgW"D��@��8���W�Q�
|xՊU^7Е�I���_�g#�2Y&60�����؏0;��yhEY�6�;<k뭷��v�i��e�]<�� )����{�-�?��F0N<�D;�#l�����S�w߷�?��fϙi�m���o��b�GM���?�.�(�w�R��D��ܦ��$�A�t���;�E����}��3ԇ?�߿A��6w��P����_~���_�̬�3�w��1��WH0
�a�h0ZV���X)�肧:d�K��X�Jj�,!�0�L�t��IT��/�ڸqCdǎ��<��~���.�l	��{��8�?�T�A}+-����ᾋ��b��+Hx�zSr��a���dH�;�Y�;���4�V��W��C���Y����@������)|�����57�(��\eŠ�x'»'������3|74���d���y�7�O�P~�#�,»��0h8��Fy�!��_�X�ګ|�"@�N��UB+4�7�!�q�M�6>���#P"��7ZY)��QD���{��}����B�T��Z�oETYQ����SN�3�<��O�h�\u�͕ � �*a��5Vs��a%r�܅.LaR����r<b�ā;��� ��B�q� ,u��6|G�~¬|��@�E��7�cQ���v҉߼-�[SI���̓�A@C�#� �CzQ$,~O���#}��8��?~ ���������������1,@X�Hƅw�p����Q��v?� ��W^}�r��~���f�����e�̨�$��`���ShǷ.���aW_}��4?����]q�,-V 1��F�(2�{o����?���2�9�9s�:����Ͼu�<����jU��G�K��	���5����V�T]k�t��u�թ]�'�ȇ��sfMw�A��P�l�CA�+m�m�޾�u��.�Ru˱"�R���ْS�Q�Qѣ�:�#�m�)��?�n�q�F֬r���ﾵO>��������ڵ�����&�F�����r� a����e�F�m����P~{�%���L�8��i���",$�k��qø��;���Rߙ4i�="�f��>�ƄZ�����B�Z�띔����	�o@��]��OvS����`Es��M�V$U�5�WB��+5�I��H��(�Ͱ�ğn��6O�|yGAbg�n��[x_��$	O�:)u�d;&tM~J�.B�Cm�j<�{�'mŲ%֥�VR_�m�n�v6{����k�&��p̐�q�Y���%�.��?�U�M�W*���&�x�����8��HA������K��۷/f���� 6��-�_�i3fd�������+�i�j��f:!K�D0�#�rf� �0�Dr��bf�L, L��0�x��0�*�5�����.<r�5=#���^	~�Yu1��?��N;�4�$p���L�?� UH�b�(����b�7������bm �� �˟�J�'�b�x"8�/❌3.���f���i���A����Dɀ�2�x!���f2ļ�aH/~�Z�pˀ�;+)�+��6m���[�h�3�̒~��>!������b�Y����#n�G%�b�;��U����~��%(Al��c�=� �}��n%��$�X!<`���c��܅�e'_AB�mY��¡�4da�9�\I�0�LDz�oG�𧮣`�&�� �jU�g��v�*k� ~t��.��'
���<�M^8��g�59m�ş�#n��e�������b��t��b�7��+~'<�pLLH[��A�c���x�T)��^{���9�����wz��.�R�L�#��� ��ܮ��_��?%�cKj2L�<���([m	�D�0��*x�����V1�@[��P�C����a�!���V��M�>I}��j���>��v����M�1de��K[���P�g3�׺uk;��slǝ�ظq��X���,�j��+VxX��!x�d�6��J�ٳ�>����}l�W�v�}�Q�k]�&��vNm�Sp�n�i�mR�*��k�����Xm�f��0l�c�F7���Ƕݶ��PP�X
�,>b����Ψ����wV���'L� �\'�`�|o����J���ӄB��w�El�h�'
J-��'Ƅk�:u��p�|�P��u��!����L�*_��Q�Z�j-�k�͟?Ů��J?�i��v�u�nݺ:_d�'�<M�J���Pi'�÷�`b%��3f��?Sz[�=��3���/�m{l�
R�N[��4��@��߯U>���ڊ�����7c�-v�'�7�����Q����_~ֱ��EA�������k0iʔ��?����~��%,��0�U��-3Lٟ��� 3�A0�W�3��|d&8SfϘE#ݢ�p���`���<5��3{�����*-ݞx�	;��c<�~l��r��U���2V��W�"�ɰ�)H~�G�q�>qH����U6�l+*H@2�j�J���N{>1~��d��{}��	��&J�N*��!Δ�[�b�.��c]������*�5�*w�m�KZA`���qE�`��@N8d<{�L[�p��E� &����Q�.�@�ls��2�3�������$ۂ��-�mFLj\p��v�q'Z�5f��p�ܩ��*�/a�uԨQvם�[q��޽�B8򦌬�'a�r�x����)G�C���y'\�����)��3����	G>Q��ނ���uy�!p"����fu+~'/���8�#�Hg���Xa ��=~������b���tķ���dQy<�:���*�N;�h{칛+����%�ܓ�,������%��Gy��m�?�d�9J�s��m۶�����G��wp`f��hGVF���ӧ��Ի��7x�`K����Ca�K� 
R�����D[M�Ϝf˖��&�;�x[�]���P�����B/ 9a�/�-�H����zS ���)�s��1v�y�ڽ���P�G�]��[���˕��s��c�=�t�b�_�1��+�(4�;��v��6�B�S�C���q( (K�!g���]k|g��J�]�.󭈥nX	�U��o�]��t�g��˯�2�R��?ˮ��
��;�_C���{�+Hq�^�A&�e%�0�?xuO8�C˴7f�)} �#5�y�����Ͽ��˗X�����Kֱ]+S�}��O���o�ci��]Ab+�z��1���įd���V`�r)H�$�Ial�F�-�Y�5�{���m�������Fa�1n9�c�?�	�̢�,@��p�ɏ�
������6~㏰R��DL�{�� ���p�Ν}��)S�w�,\XMw�/PoB��n�˓�a�/w!\�[.4%�G2�v(�����$6$qK��'߄O �G���#�OQ (�i%���@��1����^g��@o�-9���oLx�b���Aea�p���#�0��V:���� �/�1�<8L�kL#3�#�qΠ�p�5m��g�;th��H'����^�[��%� 3��ǭ����f�n^^����;IP��>�P�	���+V��Aj���w!�갅��,L�2��;��r�P�dP'��<"�pH�+�!we�����FZ!��������P�.=��'���očg�d ���Ov���K����	G��͓0�v���G]�8��k|�4)�Q��墜��R���z�-��}�W�^�L�m���s�I>��#]��v���G¢ �gQ�:;w�J�L�+1��'�Dɸo�m�f�e�p\�;B� %�3LX:�Ѱ�C��v��9������ve�3*^�ի/�9�G�t�z�� F#�:�5���0��$������x���~��&Hٚn�ǌ�7�fΘ.�r�M�8�&O��W �s�9�k0u�<��o�ǟHh[�����@��(�;��1X1arKz���PN����ͱ��Ӆ�<��|�m��7#�mނy~���5�Pdj���9s�v	}�N�	�Ej/����g�]��n]�Z��9V�nk �s�8r�1� �an����	.An߮���jڤ���1#��<����$7����֩mu��X})Tm۴�]��,������˝�qn:��/��+h� �b[/eP���MXp����W��ꗤ�~~��_�&�|�T�Ο?�0�߼U;��ìn�RMt3Y���Y���1(ƙ򱣜��665�Ơb:�r.�q�jd�+ �2s�w��w��w�-��Cy/��u8����k�ѣ��\T�$�C�U��� �0��Oh��~:�Q˅j	b*0z��b�~۳�#DF� ��Kh�?^٦����9���7oj;vӭg�4�0������f��f��om>ȇtA'>����*���!nxw��N<�;O~���?�/��O��� ������U	�����Oey�o�fy#B"����V1qU(��"D��&Y ��q��_��mI����_ɯ��C}Vt�o9��bz�4�_���N����Åw_-�����S��`�E���kܨ�5j�К4n�kӦ�-Q�M�8A���Z%��jdJ��oM$H��.��@a������\��`�6X���.����n�n�mG�$�`Ar�3�ƌc�|���"�=j��.�(���(�� Ԇ	�@��M��� �P���?
$ۘ�A���I�P���G�P�8?��Ԟ iA	��׀�?S3A>a�j��'���%�������蔚� ���=���o����>k�|���O�~����
l�$2&�9���"�����?w�����҂%0����6%��!�r��;�fHP/[�ھ�v����W����[)�Ӥ��S�^�fm_(-].A���j�FBu��բ�,�]�ǓYsf�����5{�o#C���<�UFtf���E^C�D��=C�7gb�7k��	�|X|��o��VJ�� �i�Z�s�o���{־��W����ocǌ�ys������U/#l���6��a��{�z}4k��6h)��ܨ�����fL�.���bw�a�z��oy�3����v��}������g�}�[h��W4�@�௿���G�G~do����=�~��W{���A��Ρ��L+U�'J�cՀ����c�?$�N��G�?��Sm_)!P+H���m̐�6^�g��I������{]6�>��3�����������n�w6U
%��S�N�mt��Ғ�l�^���
��.jhL�??�>�d�xV�V[��{ڞ{�~�:rC���q瞺j���F�m���\)�X"��8�
�`B��J������5R��2u�����+S�z���F�7�񃥰� E���VUƍ@��nS`S�m*��/a��a|ߩ{���֬�v��-
ҟ�(H�\p�EU'L����~�STT�Y�^}1��0+��CǓ��[}��n��.�t}.o�p�fd0�D�U:.(M\<���6�mF��Y1�`�����1s��k��z��e�7��S'[�w�y:,ջ@�6ՙ0|͕1g�>�i�
�[��'B63�@bA��� �����Ŵ����A���U
�>� �0�ӷ�=g���~DI8��rB�Wt����y&�)��w9D?\/L���t�����N��c���_p$��������gp!9�-;$�P��I���UlOҍ����U�]Jĉ�J{�vm$��2P�/�e
��3#��E?�!�g�1��:H�mצ��E���H��ٵl��iRhFy�4��5q�D7��%�s��ve��0�E��{�ys��Aj.Fdf��G�
��4c�4�j6~`Å�LFP�_(K�+���L����7���f�3�]�v��<q+�+]k�+�'$!��o�6�_��΁�7�۔��|����ah�࡞���gE\�D:��A��Ŵb>����"-�w\L'�58�������|@~�D�O��������1�Cs$����w��va�څ�ge�ULf���¥��X�㉲qXy�pV�����O��"pWϊ�WX-e�l�hOʩڸ����ծ]?����С�5n��fJ�a����eV"�"!�>��`*��x�G�l!u��c�E���-t=��=��~��x`͌0VZ[�l���٦�y��nB�e�Vv�e���{쾻����{�N;�l{ﵷ�辍��/�|�

�yM7v��A���n9�:}^�8`?�~��f* A����LJ� ���{�1ַ�~���h�|�_h�ۮ�ٮ}v�B��ڷmg�~����ͳ�E�S��.��j/Jib��93ܰ@V�l��di��omڔI�$��~֫gO[�6��P*J�/w���_�{��>��=���/�gc�H`����V���p��U��rU�X�C�!��a�;>��1}��"F6�iOH����1���5jo����Cu���'р�{Ȑ�\	KM���j˔����:⛋E��hh�����Wh�)�+�Y��Q�C��
1����.Yu���w�%�	⧃T���!yx_����	���$\e������3�AZ�S|�WVy�I�P5j�Β���o��EA��@]��f�Z�ZӦu���իV.-.����0��Yn�B�yb�~'ƪU�}o8n�J�&s�
������`�C)a	&�X�6���yX�X����&�9i£��W�j��Ω/F.�do7wY`)�jf1��(,��'X��
��1h �� ��/@��$�|��X>�+=�R���
�?�� <iǨ���ض�e�x�e���E�@H3�1q�`v�>D�n݆V+���y6c��=s��ըi��98�gJ��Qg8�JX��gk�)w��H�8�^ �aER~�S�.�:3�C�_���G�C?����@�����A\���w��
�c�b�� ��L gX8_�?�����B�g�%l��i�o� LP8�'\L�g�;LHT��K�5ɴ�÷rW��������y�ߔ!����g2�<�I��ᗜ�����x9���6��X9�nik�u�� wư�
~Lx�0�h�s�=��!�m�*@���\��n��n䀭z����ξJ��xi�cڴ���jX�Z�����DB�b˩YGJ�RL����mK�K��T/��S>��/���c��|.�h���nl`�?����/�������y�>��;�Gi�_~���N֡c{kԸ�5i�Ě�hf]��b;u�h!�5����{�|�A���&�*��6�G��{�k�?�[̣���H�?7��i+����Z�9p;�Sl�����tr��(K!`+|�-� ��k��G��F�7[`�gX�c:�rٚUR��d�G?���<������]o�.����K.���!zA
J��W]�w"�s�9^wV���k�.��O>��;�<ảO�����w��z�)R^�a?����d �
��~��T��O�����O9�Y�?|�Qq���n�
mch�Uu���ϛ7�W�xK�a+(
޾��+���+;�(��V��[޾�'��Ta��-
�f�5j�ege5I�����2w������m;�4c���&���a`��0�3bOuAA��H(Cl������� }��N�0:fv�a�<�Z5k�@ɶf�L�W_-�R+Nl�X��¬
�O�`�k��8,_1�vpF(dF�H��k�5_��w�wΠ r��
��a�8�)�@���
q��ns�'
�@2��ϊ�_t1n��H�r>�)HN?^��(�*)�%Ֆ �e��M�����r�F�����J���9�Y�֤i#	u�jXVF�[�;蠃�^��ֵ�6v衇�l9�V�X`V�-s\Ly�g�>��+!��\/7�ݮ])1�D�RT6)�_����@����e�tN}�U���j��o�m�=��o���r���P'�;�T��~I�����d������F����6"��a<~O~��:���T1-��lrT
#��X���+W��	aC� ��O �bYÍ`�#�0�t�4��*�%�\��q��:�������=�Pg���I�Z���N?��z���U�N�
��64��D�l�i�ts�����,�!{�h�zu����Ů���Rp��2�0��{i~ �[��*�AI���H�W_���K@�U�(����5��R��P��f��)�
P��o��	%�)�̈́мi�u�N��9ҷ2�78o�p�\+))��]1�1�~��m��vc���X\�J��_�^,��E,���H���6|�{��7m��Ȗ�.Ri{x+�(n�g��Ɂ��.�X�6�ſ��P5j�
94~��e�>֩cG�:x��7��������$��`�� JS���xKy�I�'����v�qNg���\�{�+�(Ϥ� e�"�� �fl����������\[i�:�����;��S��g�:Fu�VI���O:����Fa��x~b���B�H���*�Z¬��`B����_KX~��I�|� y_[�F�U��ki	֮]�z�p\#��s�<H;����5�y��My��yEG>��L#?�C<(Ee�xI����2%�B��S��jP*h?n���͘1s�E���l23�l��0�g���d������>3����>h��2`V��JP5ذ^��9�e��Gzb�άP>T�]�k�:�|�Ȅqc�^�n��F;�ӬVv����@;夓�XJJJ��Qdh��L�J��j������Č�ǃ�X.�c�<My�5�ꍸ�d+@��Y����I;,�$�Z'����-�� �_����y�[�!��T�2�acP1�y�U�	��6�CPY*ċ��Q�?���XoqpM�ϰ�+�#/���X��3B<*5 l�[P���yuԑ.4�������Ԛ5i�3���oؠ�+8�$p6k�\Bn5��t�7R�A�8�#{��\X�e���1x�')��k����"��Á���İ��9 r@��g��6�'L�%�U��m�<[�H��I'5-L ��3*0���:�7�Ob���a!�'a�
s�I�'8� Ҋm��D��.��������$��zW���b�M����yF U��L�
��Nx 9����</��'�%��#�/��'��w�rRV��^�#�Ex�h��_�gԏ9����yކ�a����C-����Z�hi5R%ܖ��@�'�t��[��+ξ-_��@D�̍�4���|�v�`߫WO�{�}�[o�'�xB�yg�^��-&�r˄�#8A?��IS&Z����޲��/@���{���v������k��^Nr&~�.]�x��ڵ��~�]�:��+4�^�w?�q��cǹ��7�x]
VkUXPdG��F�04��^�̞z�I;ᄓ�;����~�5l�
�>�����\Q����S�?�VO�0�m-$P�Q�v����l��J߀w���K�^v��y�=~n�1k��������z=��1���Z���m�����[n�I�jm�S����=�=%����J0t�����	W�/F�2�K)����}?�[[Z�D��u��F������>K�1ת�V�����n��z�^5Պ���5W_gO>��5jRO�H�_>�c|���BS�o �|�2�	},77ϕ#p��2g�y����v�eW���a͛5��^����C�����޷K.��馦x(��7������%���o*��1� ]%�Rn.
�h.�EV�Y��Ы���̣�>z����=TJ9C���t�&S�N�9cƌ]4H7@I�HYq�C��y��T�&�\U�w
���Sp�W�X#��B���[�Ƃ�%��p �����FZ�/��Q�\Y�p�['m
���)0��4<�>���~v�w}[�8�� U[������yyP�t�Pe��q�~�'�8�+�P�} O
*��RR֤���eg�T��S�n��ݻo�N6��	�b�R�1�����U�7P:z.#��w�r�F|��3z�x}�������6���~�QQ|�_���;a�����w�n^p�/Ͽ��+v�ŗ:#G���]�! ��7���c�"��Jx��;Y��]��_~������4i���TZ���L'[��a֝r���/��O?)��>k�jc�u����a��:a+B� ��&C��P�I�z�.�|�a#�b���71O�v�����7!���"��Z�>�1~��Q�**H@r��f�?i � �CC(l9��-��]�ާ��~`�a��ǞRZլYӦ^�X��������l�y��~�E�A��ާ�ɟ����q�L	[m=���3E���m�nAP��C?a�E�s}K+���P6�CӔ�Ԍ4O3�@|��,�@��	Pg����08 lQ�#X�tq����� �E?䷗A
R�|����͙��ABgY���K���?\���GÓvL+�S,S�_B�D�=8ӆ �������	�(8�&��z�R�o�ɇ�[(l�D������ �<��L�6(%��j%wV1��ZL<�Z���#Ή,YV�&��ӻ첳��!�g�e�?���j��7l">&�� `��.ǎ�[����؀��|7�=��툣����<IQD��)?w1�a�zgK[��T��N�slլ�5�MMcȂ	�q���E�o���ꨥ�*�/V��0#�w�{�|�	;�S�;�_z�e��#z�ْ~�!+Ρ����b�b�����%J w!>.�.�h6b��6l�p�e�OZ<��#~��)���'-3=(1r�M7��W�,Yl�w�p{��Ԫ�
ҽ���JI��ͼo3s�QG���L��?�	��� Wh(��A�3�Y�]�裏l��a��L�8�w^�q��v�%W(|�`y�����/\l�W���o��#�z��-Zb��{���e������@J�<��g�9�瀏�B������0w��u>���H��"/wg��!J�*���-�IS{�m�������GA��'�I�2�6���U�*��@�t鋴}%*H�=9
!>;��+�<�o߾[�?	Tha�aÆ�Q��+�x��5�Zը�ZK���}��|YTn�:
����8��S,4��L�B,('8�0k�[�� �J����3�D����~���/^�G�<�B�jy��YX l��h�ez��3c����Z�p�|���hsJ%Eʊ:�Zp3������� �G��o����h��5�]+۲2�BG���*�DPf��Y���U���A��	���ߔ�9pgP�ܘ�e`E���[������}V	�I�� 8����I���C��j����>�w�v�A��X����{l����<�R�܎�^vf�HwqQ���~���ēN����gĪW�.F��e6[8a��8_�`B�R/Y�5�sϱ>�������֯����%�%��s�����u@�ȓ��)��3VB[���ƀ����t �E�{@��6HW!�?J�"ж1��IA����p�A�!�=�A��;�腾 ��oK�����~f���ٚ�{�a��	]��J��R���yü+�\������"�m��rQ�F��+C�R�g��p�4r%e�B.o��q���2Q6����R�T��ʟ�G���B���>%-�F�T��W�&Ll�􈃋�y%��uT�1�4b{���M�\)��8D�w�Go�bX��|OB�*=�c�%��7��o1lr"��/��7W��E���W��A�d �(�{��	r�<>��?ۏh�q?
|��A! �l���|���~u90���f�٬9�\��f��R�+z9��3�^��WemU�:y�: �X�;�;���_�s��6��w�U���H����O����^��c�zn��a�~��+Z���߸qC���l�<$���O�O<�+(���~)V�5
��J�.�N<�>���$�{�����O�������7W�{Ϟ=\9`��#8vۦ�a���Plq�4^��K���#�O���Zkݦ�+C���?�^z���U��c��.E��ev�	��
翠���]w�u«��7U��Ҏ8�0��7w�\�m���bkd����/ Gd�@��jP���i�aÆ����	�]A�����K���a���⋤ �ڲ�����{�[
R���J�����q�ڠa��e��n��q�&ؽB��H#���3-3��$�hV�P�ᙄ���ئ[w�k����{�����K/� �;��z��v��Y��E>1J�������gP��D�\�v��7�+�8s����
sv�yC1�K$�(®�N��NPC��}u�*x�ʿ���fgg�R�~�*�KcIQ��M3K��������aÆ����L����ᳲ�R����oa�m�C�$>�3o�ǟN�ݺ��7�����Za>�C���q`2M�4v��kԨAJ���R(�%�\?�p�i�A��կ�a����tɃ|���5�5Q��ԭ���T�5�,��V�>�.n��Z�u�[����������p+V�p��JVy�,�N�� sb6�Y�ȴP�p�AJK��{8`.0+#:3?ghRj����㏒S�˓N:��6�͗>�ӫWo����EEK���s��͐���&����s����\@�w�uWÔl~A�M�>�۩a�z֡};�-s��_�ه�SO;�n��zۺ�V^ޯ���ƌ�r�Z��zXW�z�?���m)�.�r�En����?��ҩ4�
�&
_������>��#��x�!�]6�N�x�������0J1,��z��|@�`�w�)��ĉ�*$��A��}f��&N�dihW�L*�'P�!��?�/� �1��������lwb[+q��'()�>�R�؎7m�t��V3��ҩbի��ɑ��,���.�R��%˼\�#��BFyh�*G���I��a��o�I�'�{Lk�U%i'O.�`�����~��P�A�0���_�i������E���x�rP��@ 9,��O�o�˵�	G�� uO|V�:� ��e���!C�=���Q��D�E�FI�2Y�P'�;jL��oU�bݰ��Z��A�Ѡ�ʁS�}x8��h�����P��3�>k>��=��s�ӏ?i�?]
�z���%N�Q�X'�#�+����N<���HnXH�����2q���m�[|�N/����� c/ ��� �-�빊������:���;���>�h��`(����>b�G��//j�E@"~�����������z`�H媡�gg��#��'��!4~�D��矼>f�
g�ڪ�z�ᖞ���1���˯������6ݷ��9�" #G�f_|��5c<�P�i�� u�wd!�z�~��Op����9���3]�Zʋ	�w�Yq�O?�}2Hr���*q��i���1�'I��i˙�d"+��)8����1[<T\�'gP�S��,�mѲ��㎶���(�6{��V��>lF>�����O|�'NE�m��D[�߸������PY��x_���Ie�I���ݻ����g!��f�Z�kh�i,F�E�i��`�,���@&�fl��ð4���$t"f��ћ'��x��r��Q����;O�$}::���w�G������!KfMjH8B@Z�r�-��s�a�:�˖
�<}ϵ���-����uy��p�=>���\!���eJc����;B�ml^�[R����.��_�v-?T���;Y���}v����mZ�v�;���q���hL�J�����.y0�I~\8Ȁ��
���NO.2JtA���#���߲=q��W�����?�n�RZ���z\L�K{����߰o�a��W�K�o4�0�<��?����=�`����m��2�T�zu���=z�%�\l9b��40�v�mv֙gڙg�a'�p�<���_��>.���4QuXކ]U,ѿb}������)�����*��Lv����0�X)�/�a}�B�o��1���(#�Տ��s��c���δ�;�-I�v�i���.�����v�}�������r��v�UWٝw�)���U� �^���e6l��t�Mֿ�;~��T� �`����(L�4j�X}�����2�����H#�+
���u�,3<� @��*>	K���B�����4q�w���x�tҎ�SF�D�6H��b��Sg���K��o̺��7���@L���z�߂�G(����Շ5~���iS�y��(!�s!�;��RP_t��s!p��Y>B˜�C�E���ek��q��k��ﾶ���y��b'�N�XS����YQq���B[ZZhK�.�o��y3m��Q��;����/�뮽���/�f�լUW�l'+Y�̦N��cX����t�;g*�Y�\'�B6�T�ΘG:�c"��	�fg������˄�C��	-��XT��I.d�0�>,2�*��6ў�&X�o ze6дi3;�ē|��5�/1}��07�吒�%?/�8�4��o&[Iށ��bެ�E@vAf��_R����/�/����������IW�/ʌR�1�H��,O�v�~�PD"�'�������[�$(�����%λ��N��֩skظ��q'�(��Kk�kΞ}<h��s�]�ꫯ��&O{��ζ�n{�e�%s���vvP�L`�%������������ڏ�l�?l� �YTc�L�7.J'b��GgEHgЧ��B8�Gg�8�ҩ�Q �gV�}�0Ί3���>�@�,0��7xб�B�U�VS�*blq��mE��Y�����S���Ωc�0i�	��Zj(L�q�^휺V�����L� ���7f_�M<�ǅ=���j�V���TŭJش�[K
P]���QYQF5���R�Y5�Pצ];��e+˪U�T�
3T�UR6�dy5&��XyĽ�0uꑺ����x_��T�l�͟?�֪�`�0r�`�I���yT.s��Y)c ��@?��
w� |\��t��G�g�f�w�=��#�hF�@�l!|��g�c���;�>x�=����O>��+�@���jX���\I�2>g_=[�ܕ��s���>j}��SO>m+Vr����C��NE��)N��A��q��C�ѣ��ʝ����z�]�	��OJ����NC���[r�M���$��hJ^i&���&;ڜ�᷒!�O�d��ߔ��^���:�ơuVoX�a]�}}��x�q�+<�(l1*.^"�j���پY�n}72n�D{�������W_{�ޖ �ʫ��>l��v�=�����P�U[kҬ�ǃ��g��� ��\]��o���~��y�96o~����1[�?�ԟh+�b�K�$3+[BG=ˮY�۝�[&�F��N������#�[2��?ĥ������N��K�oҥ�?��u�'|6:�,�A�d\	q�	�^L{}��gt�Ӎ@�8 �O�%��tx��ED.�BblAń1��8���@ǒ�ҊuV�<_�"@3�V	h��~w����sŷY��o#���P�����g_�E],^z�}��׾# �x����}��Yg�a��{�a{���7_{��y�{�g���w��w�-r�����i��t��x�uv��7��\f'K18��s���JXM������ɩmo����q��`�{)3�P��>��2-���P�e%��ha�O���S�L�4Ɇ~7�W�
��##DӏSӤ�+�a[=�#�Y�q�$���U*��R�AA���\��JL	[jisp6�j]iIbuO��.;������˽R}7E�Ͻg��3o�l'�V��Mt SR�r���2�=g�p(�x�!����G}��}�U�7�[�����*���w�Q>�[ժl�GAZii5�Yͬt[�|����J��[�p�M���cl��IR��K��"���>�X�$�z��Y\��E����?����c睪���Mՙ�t��<�֨Y�Z�>�Z.eg����W�*����k��m��4��������gO<��M�8���i�����5�#�ׅ��-V�rj�H��J���+⚌��"o���	�I�|�O�'�5�؀닀Vj�,\�l�2:
��0k��ƙav(�a¡L%W���1��h	�4x��|���I<H��~E��(H(:\�ǽ<\]�L=�̑R�%n�Ixΰ�LO���P>(;(8Rv��ϨD�E�`�!!����!l~s���U"|�"���JOUgBeR�{,M��U� ��Y��jJk��V�x�o�X.�����o�Ǳ���\���9K	@�%��ŕ��Nr��PJ��e+��+Ō�>����z��i+���q��\i�҈3xl�++ے8�ʅt+�F]�z��1m�n~�ǅ֠w^�v�;���' .��eW,-��R�ܪ��e��6)bנ����t�K6�Ι��HX%&�J���#���T�6:�:��>T3��x��SiA�O�|xKx��\�|`�7`]1�"�����߼�L+Q"]�}`��� t"�J}R����� "zcjA�"wl!�1)�L�^��53�����b�w��L�ԭ��4ld�[����X���� I0S�NK�]gYzFM��s �+�X�'���ǄH�:TUR"�H�h��B8[�X%���-,������b�iO�_����wpQ��t�_8L��j�K�1~�/I�/��?�!9}�����"n��g��$�����.��x���G� ҈�q��x���'�F��T�VU��FaU=BѢ���q�"���KL_D�.<۩#�dl�f��7A<S�x?��26A�lcrԨ1~����ζ�;ގ��׎�����{� ��ڴhn��w�z����ۻ���k��l�KY���-{��;R�^��y�^}�5{o�������Ͽ���Xs��".Hf��m�L�͟;�f͘�n�����.�hj��(��@��R�ðJù,� ����{�]��믭XcF3�!>�Z��NNM?�b�0I�	|���x"��e��n�o��6k������k��� �-��j�@���w`�c�����iSmĈ���`���V����)�2���$��q��9k�$+Z���Mޢ\�3w��5.\��r��`���#P#�W��P�T׫E��W�^kܰ��*L��"���]�Z9�*�������6o�lￌ�S�b�p��'ۉ/.2!5k�������1�bܙJ�p����B��ͤ-�*u�z+�f;��ŗ�������Q�nD"[2Lzj�5�"Ԧu{�y��l�]��^=w�&����%6����^�����~��J�Q����Y>�^#n����4m�I	o��Kx����6<�t�	'T�8qbNAAA�ŋ��Ѭ�_����jڴi����ϝ={v��.Z�hi~~~Qaaa�����-�s��r�_��+�͛�\|��-S��8���5k֪3f����
�J~���N����������W��S��eJ{uqqq��5���o���Z����K�,Y����,~�6y̝;��$m�'wa��ZCx����Z�AIX���4SԩI3e���|wE@�k����]�p-gT�����(2���R��N� �����^7�ӥ%b(M(?�|F�m<\<fȃ:$
��t�E�E�\��f��C�F���V�`޾2&�F�<�rl�c�<g�zt�a�srl��I���YNfJ�2�(o���~�QGj0��G�6�>JXk�:��Z�Z�ʳ���d��;425�R�_|��}��\nչ��֧��瞶Ͼ��ߙ3�IA��2�Y0�(�����6�y����d�'�� ~1`&�y�'���aS�l�K��>��a�}�`U\�I��X� Ƭ3�I�'�p���ɇ�<�9���'h5⇐W�VM�=�s������{���P�{X����`Qc"�C��r�=(�Y�7�UX�&ҋ�\�C��YR�6�p�3F�>�R>p".i��ȗ�8��k(Sت�.O�.����#x������@,o����[�C�%ߘ7�"n��d�q�y�� ���w�G�Hg�i�'���N	�NT?!<�_��2�$+.<�8Kڹ�V�߾����+���yq���	��'~sηG�����b��ek�u��ܠmժ�ڤ�Sla�"��cKu�ڵ-+��h��t��o4V;�rᵖx4B0V����u
�:����2���~(͚7������:�����Y>Az衇��8�ӳ=�{���3;ت������Gpb�QYy~X��������={l-'=��{�Q֮m'ϛI�w����L��z�ֺE�x�I�����&Nku��1�5�lЌ�T�~��ͪר�g0VBy�z�:b����3�@m�U筥`6������K??��̈́^�v�쨣������"|绕��°��}���V���_F������n�:������)Ik9��}Q���`13##�����/�s]l��c�Vm���)S���kyYƍ-�Yi{ｇo�t"���1�C7�����{X5�lY�}��6f�oj�t�q���>PfQ�Z�h�1["�~û��Q#Mu΄7o�,Tj��i3�*�c���զJ�*,X쓭\�p�1G�x�w���>��8��/�>�_Xt�6�OtB�ľ���^�Tߙջ���Ζ3H�@Az�7J�?����h#�
$��K@��At��ڰ]w��Y	�rrr��]����5�B�o��}.����OYYY?��Gggg�(F��~�T��S�5(���x�f����o?ԩSg����QOR�q�6Z�F�}N��*�(�3J�1��N����w�S�c��x��;i�דt~��	��8&�N�;���9F�ؘ��&��D��K�u�i�L�Jo��MQ���9���PL���-�c��&(����0��{��9L��o��=[�i���P]�默E�Ϫ��<(*k�$7���q���g��=�+3�͡����=�jљ�#KX�{b�j^�D�wVpTK���c[�s�=��9���gd|�:����n���#��s�o�F���>�t�w�U��p��\$F�X��1�R�U+�C���~f	���i��K>�g8���0rf�U�>( ��@�Q���K@eL��Hf�t�%�~$`���3*H�����M�
�� /���7�쁾����!,��vq����:���ąN�AV ���ŀ� �4�z@���H|�"	+$�!̑N���;}��0�X�<��Hñ,���zR��o����o !:(Ai
����or���ő�	�e3�A�On���3/�!n�o�31��ؘ6�yGY"]��#��G����6��2.���ƴa���w��
@�1,~�G\p@�01.e��MN����	e	8{=)l�#���#|(K�Wv��`.6�"����R�^�����ڭ�1IFGZ&uM;���2�%�ij۰u��6��ގLJ�ʪֵk�Z�)�5XM��Qr�k�+|r |)3��w���ğ'8Q^Ɯ�-�X�c���Ύ���� x���^={�Ǉ���v��=�8���6t�P�cBp�6�'Ǹ���G\�p�|;f�x�4���гgo)ڐ!���J���8)L=oƒ~�H)�h�w���3����R�&���k�l�U��L�={��R.�j\tʇ�~��ER6���9s���h�թ�@���ו��ek�����Tl��jcG}���� M�>�>��C)1*H����53�f?7��8&��^���f�Q,�����:pfU�6FHKϰ\ѡ+HR���w/�q��St-�6��x�GnY�ե]��d{쾻�kU��k�o��#����<�\�ee���'���]u�zkӦ���nůe��ּY�[#Y|B�C���0l��o��N�Q�n}�m�(?ι룎>B�N���j:�{W<#��7���ir3S������?�q ~�r���k�-F�D��5~�ؚ����U�Ұ�C�%"�"	֫�//��#���� D U5(U1s�Ɨ�*z��G
ÝEP�_��w��]��G�t���{���)���m���`�,�q��%-\",i��Z1n�SIx�MB�_\+��4�IE��$�r�08$��*R��x3x�rP&��I��V�/���	'�N�T�OU8��VW��n��;������^a�;f�+�g5�&6���3{S�j��s�3���|g��ʀM|L2h4�@�>�)��{�Q����b�	[/��	<������:SyOC.�K.�Į���)�wޱ��:Ƿ)����Az��v�!���/�du����kv�y��*[�k�"m�}��Uv̱}����3G'O��O9�~����:��Q��j���{ہhmZ����~�.��B�#ISn���?���$ɂh�!P��o�I����K5~$ A?� �(E�2e���(��R���� ��6��[2h+�_As<q(��1,@�b<o��r�md��3�J�#3+C�Y�Ҭ�B}|�7���$���_0��� �"�h��P����~�AX�ȏ߼���x�I�L����I���7+[�*���C��-5p��+<�I\[�%e'?�g�$�O�Cp���'�\�Vm�	'���<��uFx�!o��tx�e�.���>��	�3��7�G|q�v���� M@ڤK���� ?�p��6q ʉa�㷯b�p1��KߞW�ɚ�,��!ps��.;����zǷ>!ܣ q��/��;P�Q��Y.���-��A�f�J��[Ӹ��M��˄J*�*lyCQr�Q%`u���jU�c�$�r�-��RN� _�c]�:��<�w��8{إO/��� 	�M�>�ڱ��C��̭�a!rIq����s�}λ�}��4��^׉��N��Q :��u��GI8��;M�r�I*S���^�{�`ziq���{�}�� �]�k5�=/�a��ߋ
��I'�a���y�ɪ�j�����ֵk7���M�0�j��t�:O�>�����B��z�s��O����a?Z�~�ڒ�|;��]��W߲ZY�s�}��0;��sl��1��ig�f�<�e����x�	��oW[���m�]\��m;�a�]|��x����2eP�y뒥���r:�;�\�\��x���ŅKD�#�_�7T��v�=��e��Ua�'DOO=��]s��ly��?�������(��Lc��n�&-=Ųk�[�����;n�޽�(�����xK_�'�7����!���^�~��';�̳m��_��_|�W;Q ����[nv�-(�o�'���f��]@~���a�<�~飼�%��񞑑1���?��O�b��O��t�ܥ���۷��3>���:t*@9�[ZZƚ��Z���22��$��\��%t�k׮�8'�NA�:���֭��{͚9�r�-�W�A�����/�0y���S���[�GX=��@����	�@i�oРѼ���ߨQ��J{^��f�͑��G^͛��ײek��'����?ᴐxM�4#�y*�<}�Ӵi�b��6l8�~��3�����5j4M��իWoz�:ug�,s�����ʪ������`����o�c��n��}�N��/��4s�\��]_}��}��1�A�����Ïr�L�ε�cƸ��3f�Ikg,8��d�G����0��h�C�A:y�=
��% �`@ ş�#�3�E`�X�IfW���g~�����˯��n��}��|V�!`��i6{�l��vv��g��;C��/h���3Z�j�[�a�	$�0��(s,�?1��*�U���d� b:���\���߫���$��$��$BҎ��2��?�/�7��;������h[~���I�H���6$���WL���R��I҇.�'�c�;[p�ρr���:��'�̀�� ���<��#��P~j(>@>��!lA���]w��[lv�i'+� W\���	E�Y^��;e"�X6�u���Xf~s� 
u�d	O���ń	
۾Xو�!l��l��1�ے���tp�QV��w����n���x����!����H#��<T�X'(~<q1m��3��8'����4	��O|�\�"�0cN�._�܅k��Zm pS�+uܾC?������0�]ۊ���2�|)ќ]�*~8q�	�����'L�����{���6i�D�5g�͝?˦Ϝl����m�l_��0��<�;��:�>����\-�i�	`2�� a�1`�.]���2�w�x�RRβ�N?�N>�T7hr�I'�1�k�<���#��}��߯�`���p�B�oE���y��9�G�ҶL�'yF��}�-[��ۨ�l;�+��q��kO�;�Z�nc��vp�~����`ݺm�6�E��6�U�j�.>)ö7�R:`���I��� ��z G�%�������k�hn��a����k�����s��6RySE?+}r1���o��؎�J"�P*Yq�-%�{=�*FN�qL������Wh>�DHAL(65�W��Lx[��`'+k��0�mh�圖3��NV���$�
Tpk�2!����h��?�L>О ��w�+�f#���!�����6�ק��-���ol���Y�1�<�ȼ���w�qv�1�Z߾��I'��wT\rɥ~���?b��z�]q�_��/�����M?����֛oـ��K/�dO=��=�����7�|cc�H1@0����g����"�-oaۏ�.���*��y�n���1D%
��.�S�v����&{��쩧��O�>��mi\�̛k���Ϟ�<�MS�o���]�~h��s��m
�����C�n�5b���ޚ������w-$�Ŀ�l��?�Xv�C��A�A��1�1�eV�W,v���7��{[�<�(�����Ƹ8��U���z{�g�矷_z����o�޽{���L:� Ξ1��̚�P�('����٢�<~Z�h��X�[�fϜaӧO���Y�f�yBp'��v�;>I��{|#<�V�;��Q���(E�{�6���
��#apģ��-
o"�.�N�97���#@r9*BE��3�Ƕ��� �4@���xP�{��� qb���T�<����:��dx��!�����"���g�����V5�Y0h�{z^z�%������w޲����uhc�̱����}8<�Ŏ8����슿^a�{��p�	��.�~̱G����!����/�ٱRD:u�d��6{�los����-����L[GH�
|#�x(���`��z���W_}��}�]?�������&��d�'N�����̳%\���u�����kl��qB?4�v%�4�"�_2�Q�(��J�ځ��c���L�쫧��}΅R�α�O9�N9�,)n��qǟb���T��v���j,>�N?�t?_�A�zRd����(�'�	���껒�}�U*��V ����O�>
nLBGi�\p��~�Dyr@KW�P�Z�l�1%϶b�Ͳ��pۋWmݭ����u�'y-+ŨF5� eg�d �ա	���CU��;d�P������6�(Y��V�mϹ�Z[͙M�?ΕE��G���ľ�+8�O��@wq�yT�/���k�[��[��$D�),��/Xˬ��"իo�5��$g�b�����m0P.l�U�������0��`������J�Y�ԙPuuR7�`��;�1����� $�E�d�t��2�a��1�" �2/!@F�����>{٩'�`�۶�jJsμ�v��w��/�����٤k���^z�e�I�jP�'��r�����/��f����@[m��� ��:ZH�o.�\^O�N��B���3�X�C!`��G����a��! l��C�C<��� �ň�$p��~�<��dǟp����.� |23�(L�O�8�ͅ������n�ٙ�4rΜ��m���~�J�X���X���/~���c<�e��ww�����e,pn�o��`NݡDQGQP!O��|�/���F=��7��;�E��iD�7.�Q���.��\�b��U.��0��9~��7�	K�����ӎ�@��ؒE�Q��/
����V�'O�2�K+(����g̰/���uv�7���{衇�K.��1�G{�={�^`�^�]q�����s/<g���g/����y�]�w�#R��y�Y{镗�9)�Ͻ��;��K.�[n�YJ���{֎�{�ƏT7��L�b{��E��<�����+�E�<�:�ވ��x�;��W_uUb2�X;����r���������w��ە����6{V�M�aVCPJP�PF V*�d��q���)S&{���~�ͮ��Z��x��瞗{�^~�%{Ec��}�i���o؛������~�;n��Wv0�\̸�������LNFrM���X!D	��12CY1�Mv��ٺw�!���W�v�i_�b��~�Ŭ����Q_rC��<}h�'����ē~�UN)5j(�a}	�'!W����_=���0\@}��f�#��j��>E�C��Y��:N8��J�� �`{~ȑ4���%"�����	��yF�}Y�zM�ha�.�X�j��Gp��7�2d��?��S�f͚� �p��:�Dp�L�e[�a[[��ؠ �o,�3k��38K@���q� <��ԯ�c@��ؽӋa��&���A.����24q�d_��	3h�4�ث��5m�{�����d��R�1�6{��l7k�3v����Jһ���Ll��l��2	sl�����u�Amذ���[o���7�|+���6\�	HʺQ�$ֵ�@��Nl$�+��A����!%�qr�U������~$����I<#İg�T��Xn�NEp`�E`e�Al�m���m��F��j��OmԨѾ���Čjޢ<߆Ė���"_�E�EPA�B��O��y���駟"e��_�fm��W�|���Ա�v�!�p��~{;��S\ ޮ�vַ�թms�'�HɌ-�P�T�6q�zRٓۈp���	��>͊�����`e�Q�B0;N_e�|H?�x�~�R��=
���� ��jN�@�i���b~8�ɋ���M����=�%>.�I���w�#�Q����ӫ�Ea�	nn�Am���X�[������7�|��w�s��H,����ӕ邂|�4i�+�}����{챇_��4e��К1k�ʳڎ8�kբ�oEx�;�-�]h,r:.Z\�w+����� �@x��ѦM�ᦾ�r�P�yi_U��mO}P�eK�ch
�]��Rf�U�����W_yU}��i3�l7;�������^|�fΞc���qz��`��"��%K��G}��3��g�qc@s�γb};�Ŀ�v7&�8��>Rc[6��~�L�^u��\�G�:j��q[%����>��S�يeˬc��R��"�/���}���մ�~,�g����H����>����}�?�i�������Rf���M[(�W~��Z[im�7��?�2�Y�	V���+�%��ݳgO�g�}|,�^���?��~��9�R�W�ƍJ���5p�������z���g,P�-��Ol��V�3Jϑ��3�7l����Çy�쳗��~G}K���B�;+�e6n�?c��n{�V]�y��/�����kҸ��2nKY�s���;�^�9R_P��������&h|�T}ZB���V�I�4�7~�����R���J��ѯ���O;�E%
 ]�iQ��y����P1Oa!|B���(��j�.��;��[���y`�Qk��Ag��pԝ�)�Ka������H�&;]�PG\��0"�Z�x�	�w-�Y]Ÿ�I��������hʅ�fw�	�T}��� �yb��f�)C�v�=��_h��z��9�����ν�NC<��S��O�SN>�.��R�߯�ʕ"娑�V��̚6G�u��賉��s�]��k�o�\gO<��}?�{)�X{
�A1�ά�j}�>D���mA@����/���Ut��תm��a�$�)�Zz=���_�J�ʻ"���y9}�o}'jq��a0�>��Ji'9�+��,��r�'�Aw�0�F.|�/����g�uh�����=(Y���8Ԝ%�b���>}���A�l�Z�3AK���'�?��^~�>�d��,��NR����]�X�fM��dH�,��$|�6�g[V�Ty���͚X�.��m�V�ϰC<؎=��v�a.3�ڽ{w;��3���v%���!�'mPMB�Ϻ*]~S	��A�W�W��T#���^��ϵ�c��6>�1�1��ϒ[�thW�U�-����HV ����X�v�|�� �%5�&V�/H_�"F ]\���P���b����<Y��_���:euk`�sR��D|��#�������?�p���z@�C�	P9~��D"�&;�/�ёRb|�vх����_k/���=��C����=bW\~��v������ٝw��V׸p�
mT,:�vE����M���a���/��|	ɢx	�+헑?ٻ��ه��+�?��=��#���O�����-�f�7�`^��;^���֯_??���~�����ĶB�fp��v�����l_}��O=����Ƭ1���QPl��~��~Y��B���&e��v=�s���~���Ty�IIl���T�:X�z��O0v�V.O��.�P�x�,QX��ڠD3D�b浫�#� �^��G������ֺMk'�XYB�e�4�B�pˬ��,#��+d�4&�Α���q��?�C�����#p�kq���[��T�J|�U`��_������/�PX��� {�٧����:��ҿ��]i��v���b�=�O��:����`�C=�|�V�,�+��1��V��~�m���c����U�T��S�J�&�4���Fۈ?x�B��.7���; �'���3,+=��V��D��ڝ4K��DJʪ�$02�-*��9���/\(a��d&wc�b_���?$��WAEh/L�O�[P����*vʱ����63P����$1Do�Eb��[�F�K�.D��g`��F`$tPf�y�[.����`p�
wg�̧Pd2��,�s���UF1B��@��H�(y����R�v]@�|�/'��5h�X�:T�Z��`����R�p�$mب���tؗ.S�Y�3X˱��(.��2�v=�S��~g:Cb;a�ʑ��R���A���q$�ǎ����y �ޤ4#�^@P�u�p!lRJ�%� ���C�� �r��OL-��>@g�B�(�l�p]Cb�'V��)�2 ,��(H3q�B�cń�!C����F��p)I�]��}A��}�<��#Xp�'3������e�r3�����b�l�q~p����MVK�m�֭�a��6a�8{g�;�v��m���:�] ��ׄ	|���`e�"п�1���G�����eh�����.Q݀{T��Zѽ�2c���1�;p��Q���4�HO��͊gbk���y@l/�}��Q� � @�L�r3�"��3�!mA[�v���yc���H�)�d�ڼܕ�p�L[���"E���Ә��K.�UtG(��/[چ���H�{kz��Κ�hn��˖r�*�*�t1b��VR�T
rk�SV`&O�h�����vۭv�=w�g�}n���������~�=�٫��f����=��3~�j)����YY.��;S�'��r��XzZ���-u����ϹT�y�?�¬=+��31����d,�̚�|S[�N�9u�_�)��7y���u˭��?��L�����g{�k{��7�����Kh	�'@h�$� )�:	$��K���q���������V��$����G�˳��}�ёF��hFI����O<aW^�C�mk�V��'�iG}���_�!0�O?�'��@o�9��a83���C}3 �MIm%-M|�ޔ��Ł���`��r�q�ƕ����?��J;�o��G�[d�'���s~`��`��
���x�@[�u�-2R�kuE�&�^&����Ì#/������W����=�W{����^�ٳ�޾���'0@��Ass��3.<���x������f�d���O?����U����v�W�i��i�>����Ol���I<�z����ZVp�O�BmC�]�7�D�[Z�L�E�� GА�\�d�]z���_b߿�b�W=�:O�w����$����
��Oa���"}Mm
�1�D���_A_+�_HJN�V#r	��@���A����7���!��/v�<C��@!��9���{�⺇���؅+č��̈́gB��������Ý|p��?�����#�<�=�Kz�>puW����M����2˫h�1�_q��A��~��h���Fٹ���ˠW�?�7H䑾r���N-���8���6H[V�%�V:�T Jy�|��J�+
<�o ^���pJxO����-SAA��Ǡ���s�{R8�dZ���V�_j�U��nm���C�$x�D��.I,���Qx����7!o�1bϖެ;aA>�qqV�)_lc�h�B}��!觷���9h���	@v�c�Ŗv�����ӶdlRů��L�G�D���'k�G~��{�Ӟc���e�3? �c��;Ȅ0B�1���t�&B�c}^���{ ���w�]��=�wbZ�hN��z#@S}��K�ٽ�U�i��u�b�27�9���O>vC���?�i��lf����f�v�eٲ���5�c�����h��8b����1�vfP�q�Ej��+-�!���0ʑ�Q+�k�<pet�##0ֹ�츢r�l�&�(�(+<�� �e��u���4c<Zh�1CF=1�WYY�k��������S�]r��v�u�۰aC����]w���V�s�,���&�� �J�gՄB���3]j*ʸbaH��^`aBiJ�Z�2�œO>��;�\w�eM�_���p�	~��,瘁GQQ�n8��[/~��&IS���|����h�_�#|h���n��]v�o0����g��n��v�1�#߉�n�/y7��z��]=��3�o�ÜQ��<��|��g���t�U�+�wC�n[�'�j2Ѓ������'�����ڴ�������|�Mv�����0hy1���.�ڀ��¦M�ˠ��l��456VTT�H��4@� B@�z4^T����e|�"���֡8��b ���{0��Q{qTl˕�(�vY���B@���b^��q�>tJ�7
r:"#�Q�8�ϸ��8�+���w����%D�R&�"�b�J^�s�@�|\)���9|ߍ��wK� 0W��jk��[�ٗC0 PP��M��\	 �1�3"�Ca������=�49;E��Y~S��:=�M,�jj��7ޱ�^|���Q8`�C�:� _c�:�G�����p����"��a+h�]�"�7��"�O��b|)N�%F�d5��B?~ӮP|�!x�n�+��.čyF:G>�X.K���r�wb�>k��0@B������|v���B,[L�|9H�k���0 ���1�Đ��i�?x2]�=^���Q���+��o�.���� �>�� ����/��Q#G��a�lP�P��ҒVUY+c{��i���[}��uU�d�r�%y���<�%�1Z�|�
��!�>@տ��0n��	�����(e�|�n��҃u)lD����P�	2c���q���3�E�o���{�=w������.��bfp�W�W���X�x]%�$>������ɟr�x��z;:(ߢ���NR�1$|6f�?~�|P��|�m_���_v���/�'p��Ó!���CQ�2s+�7j3�<�{�������!c�Y �1�MY�h{�7�at衇ڥ�^j촹�;��{�m��~�� ����z�=��#P���c� ���"xoꔩ>�����Ķ�e���b<��7� ��x6/ ~��Æ�*c�h�m�����w�6σD�o��?$��M�5��?��`�����ς��C�}�M?E��04@"/#L���bD�PB�|�)ݙ�\�q�"�*�����Qq�~����A�d3Z���XCP"X�7�8:�����O��vޣhDE����Y�qb��#��1��&D���!�������A�ҡo,��r@�X��h�	AU��6�Mb������-�GQ����.(���1͘>JP"�B3�aCZr�rz��ɀg�Eek��%nР͝3�f͚c�-Sy�l��aR G۴�[���R<_}�u?����C��]v��&M��ϟv�i�����=F≏s���7�ǥ�uGS�L�ݧ0�B9���_�@��N�X^B��K�c=C'6z�nS���č�Yh#8������f� �H�(�� ��j_�8|ϻXo�s�8{:���w �'o����'��K����yĐ�/H|�@*<��B�;M�lB/~3;��P��~�+r%�u���y���o������`@��x���s�If�Ǝo��M�rL�݃n�lV�Ng��E�c����8O����G��{�1vrCI~��'����+�}��2|�v��<>�_�̷�����y������ɀ���2���cF���Ϸ�o�ݶ�~���r�1���) ����t�����dx/����5�jG������AE8\���_����ы.��n���j�Ci�>�L=0�-�Y�f�����>����v���X;�#ZYt�B�����=x	��:c� 7ؼ�g��5���կ�؁|Ў=�X��� ��h��#=� Ҡ~��B�=M�mA�/!,��m+��!ۨ����������>�F��6���^��m�;�m��ܠ
�v��/�P{��k��~Q]]]vgGG
B������0��J+
&�0�dB0���+ۀr�(�&�3�&O��@�^�p�1.��A�����9c��ai�=��&�!��"o��{��F����x�G�ߠ$
�(Px�}��M�8E�J��;���EH̟�I�k�.�'��3H�y}�ގ�{�%N�0���d��8�ni���ٗC([bHL����� y6,g����y�1]`}��&�?�	p�/��m��qQc��0Љ��]"?E�I��ĥs�}9�7�"0R�B�� ��`��� .Y���X��Y�6m�r����� ��\����p���>{�A��켫�&�v�6(*(���!���.3V�﷿M;���f[7�hC\i{����	�|i�rx��ې����=�󕖖��(�>�%�''7�

93�����0p�@+Q�R
�]
�z�&���/�3����̳�vq�\	�n��Gb�X����b^���;��
�-�G�+��r$�%~𜸄��oQbI�Q
�(���C�g�g����'C�>d��j�=�~۱3���
���O<�g/F��5�$�.6�|�3r����^{�wl=�y�A1x^�9���;�<��8���EE�-�g�?�������������#
5e%?�xC���d]xᅾ�uήx���[n�w�y��x�7�1@�����.>��g�j��q	��I�L`���1S [o76ֹc��B��3˅�1���E��.����_��R�dKt?�����W�k�.������-(����6~iko���Z�KƘ�N��E�E����]N�̬�U�Z�=W�#�v�Ln��w�{A�0�}�[2r$�k��4�W�5��b�[l�>&?�{�!����]{W��'Q6�޹�/��9�}�o���z�
n�|O�Qp���,�U}���Iy���Q�K����8��Oz���;���8}�?�7�x+C"��N�g�};*AHIx�Qv�=B��]�
4��i��q���?:��Q�x��B ��.n�˳��ٙ��P:���6i~����]��M�xr�aA}��(DH���;�'B���#������_M��D���� �!@�<_�!*E��)�D\�xӥO�i��U|��/x��!|9Ĳ�� ����C���64��y��x�a9I+�%^����f��ȟ����"��P�ÿ���V�|חo��6W.0Lv�mW��7�*?����뮵�~x�����#�w��&Naesl�)#�ȣ������|ʉRH���w�}����-{���ܰW^yŞ|�I{��w}��e���_��1��.{�����{�o��~�s���f�=��/���C�"�� oĲ�Z��G;���ٝ�v�<A��~"��������e�Y ��S�L3�&!�	]�Z��,��,�w������B�����x����#�k|F�D<�7�ac��}���o�;�.�@�������no��\������K��[m�O�#���7�gw9��G�N�j�o��m�=w�C���6u�d�j�-l����řW�ش-���������+q<��[�nl�?΍rf����j��+|���C�Y	�'f���2��Qߔ��I(��ʜYSpfM�@|�c�0B�Ӧm�;豣�I�:I��47V�w�9���=���1c��ڼpf���� �EP�kk�ҮsC�����w ��U���!Ϋ2��Ej���~��ag�}��~�~`4��_�v��ת��0���Y�*E�����=hͮx�rs�ڐ1���c�EŖ�B 
4|f�(t�F�(�)�^�� &}���Go��1���׿��������?� �A	!Cb�U��ϴdF� bۆ�#/BO�h�D�8����r�MI�+iz��@`}"���`X��Il��N��������[���>ʠM��A��_8��C�$̶�N��΄���n	��}5
HT&c`$S"D! �;܆>���\+V�(%q�! ��b+W����{=��l��x�b���6g�l)���h'0O���ǟ���:�(�6�Ǘ�w �'
�#`BtËqy�o�(F������:��47���7��4�dH�Kq��{}QA��}�/B|����>�,�^�H� ���w\�'�7g&�3�`��[}' (u�ކ�F�&��B�#���3�����N���1M��2FZ��I��@�����ǳ��unȰ悑���~������-6�~�%V$����ʂ�\�ʖ�M=!u/�X���J~C��}_����O=m��_�^rE�6E[�����k~�
�5�����3��+/���YԌR�Pψv�'��#�C'v��e�t�4 x��:��6i/o��.)z(�|�)F�雟0�)���ٍ,z���'�:��C6'�<^#��A�6
}qA?��\Bx�J�U���]�%@�"�.�=�������j�2��}��}�����#w�y��I����>sZ��8��O6K�������3<�l*r� ��Q�Ț�e��C�����fYQq��a��;l��c�Ł6r�H=j�
7�e���� �&Ͽ�}��{���鳇���M��s �h�	�+�� 8�6�r2C{��;?a���~��s�8�>���>T��"G*ξJk��]��+�G����	c|fm�ʵ>����N;�P9F:^J���ՆK�\�W��6�v�q'��;��}�	+�q��!�`���~VU]i=�ʛ���n���&?��3���Nf�5���l��v��[��m�ɓ'������D��VqU?�ȣ�΀�_x�|�ǋA�]��cw�����;]>��Nkj��Ύ:�hkk�����x��k�����hK��G�}��4�����z�>q�dM|J��`\��5x��L9Q�P�ȳ��4�u�����m��{�;�}�Oܒ1S��j{���V���R:�l&��㌩�>��
eP1[geY���E���ucm0��1�'ac��e�=�q�Yii��w��ɻ�{�9H�%��@�����R]U5���ezAAA���I�'L�
h���SN���y����1��D0�q�;�K��̂�`�5�Y�gI�pw ��~��\�&H�|�p��oFĂ��eH��l���k��߬:kq�҆0�Jʎ�����x��\(s��}!��w�7#�н/�.!
v�ا�Q�@�W��/�!\� P._�!��6�����(eܺ�<t�4��	FN/��RϹ�p��c%\1Z�>B>�9и/^��-�sP��|C>1e���E!���2���g$)�h8�2$Ҍ+��3 ��������nU|�!�x�"{H�CUu�o�N
�45ZvN��U7+'j�g0-YhoΔ!�̓��G�;���;ﴳm����0���v������g�ˀ���R���V�M���Å�5��B��*�M<������4	4�w�F� �]���I��p�-.h��Uz�#���.��{��LyA��i��ΌA���c����G���;1��_��_N'�݇��D\���F��#1@��e-~�wo�	�e�߭��x��Ј@�=�n���v�%��ޯ~}����m��)缠�3��u���H���^	F�9_�
�R�n<�6���$�HK��ٍ0/?��(��C�e$��<�{���O��3{���l��%R���_�~��q��'/��_lWap(�����_��>_}ig�q��_}!�}��w��{��a�]|�%R�?��o�A��َ;�d�z����>K���;��ؑ6{��i�%�٣U��K�%ۻ�~��5�������Xl�Gm���/�A��t�M�ٞdÆ�u��|P�~ġ��=��ÎwkK��3���v��F������~*cm��gE;�,4$Γ��M;_�j����lV[���[o���.��Cmi��j�->��ׇ��d$0[���#�VHn��1�p�m��w�}�^$�U<8���#	�L�ͮ�����+ xu���ð+m�����{v��ͭ��M7���cƌ�*�v惷��g��ߴ#���i��-����f�]0��:{����׋�A	�� ���o���gYSK�=��3��g��(/u��g�G��|Oٹ����6�y�I�X���	\$?3�_�F�THO�y睛����r�&�_��}���{�������t�&=u�m�C�>����{l�4�0�BG+��	��[�)�7�=��x��NII��e�w�V:�U�V���/�u��o�t����?�Ң�c�cO<i�w�����$�(�"�����Q�?ǫ'(E�终kL��,AM��%��(���ѭ�!��X�kb���"�e�O��o)������0m�/�� ���������N%�_ļ"�~�
e}��R��C���AaL_�*ΤӛR����_]�o=u�{����)�4y�I� ���d�5�24yE���p�S$~<S�C=�U
�t�P$��Pbq��%�'���c�6Az���l.\�ƨF]kk	�:x��V[M��S�pW4MW��}�]�zyΜ�AQH�p7S�l��6l�H+-)��F�@x��7]�j�]7���ЫCJ �7x5EF!;f��,�/�D��f)�W�#X���.���*��Љ{ E��oh{,Lokk�ή0��a�"ch�16d��W�r���M
%�]���x]��`$�	�xU�B8+�A M��7�տ�O���S�����^AfEY�/��3�����,���Pvp��H���/R6�~B�yT�c���r�ιW<��.���v�� 8���؍7��ݘX��L���}Ch4�|��4r.up���ٞ{���8"���_P��w;���ħ��r�z�� 4��퀚�Z�t����Y�F������A�х-�Y��z�+�{;'h���Q��� �0�岽t���6o�,�=�~��ۤ�?�FJ>�0�������ڹ��u8|�W�1���Vq%[�r��[�֮�������{�V{:�XK���ʕ��xd���<h�eg���R7قE�dXrȭ����l.{i�f�J�6}���{�ߏ<�X���#�2N��No� u�����{��uC���{���ˈ9�Ϫb���u�6l���q�&��3Ԙ��/]�|��av��T?<7��m�l�%K��2`1j�):��<=h�K&����a(�:�*����7�8��#��'�=��SO=)C����7���lMA~�8�����<���'}n9��©�vg�
�FoC5������W_a�<�Ʉ�ƻ��-�$Fkjj�ʵU֭�=MF� ��J�p9J��Pe���\c�9�L{��l��1��i�-��f���֤zl�:�� o�6h�m2ʉ��?K�v�Ls��^�A�c|�^ByT'�]xᅧ���sz?�_s��q�&�_�G�|���+��w������?�SO<n&N�µ�}������E�#6�`8�h�$�z}~�xeE?{�rʷޠ���\q��8a�����6o�\)	]�Y�lg�du5v����Ϳ�ن�q\}�	;���Cm` ��K(1�+	@j�_L��}��<aɁ�(ˣF��1cG��T_��t(!���A�F��`)��<'���_��3���f����R��Չ���^4sC�|ٲ�VY�8414�P�X��nvJ��N:<��[Ҧ,̬4ԷZUE��a��Ά��C.oR��3W�U��tEN�:�3���P�)��;��T��r{|7X����'|�@g	��CO"�+}�P:(�(�A�3;z�.b���M�wC^8�����d$��\��Xo��u�~Ў��鐡Cl��5k��3��;�	��'���h�5��E��̙ozG��B|F���ZfRq'Z�l��o����7�
faP�����`����x�[����RO��1�x������w�w7�\)���В ]������c|x����DxE������FՇ�t�hJ��_\�p��o����cY�a�5#�~}O>���(������<�|�a�g��3���t h�o���xo��3
2|���;�IQۡ���8�w�Ʀ�O�]h�?%%�S�2�<�%�!ʌ�%�6����y�_`7\�3�G
���n�ﱇ���}��N�!����YSC�ʺ��/��v�a{��96x ���^{�
׺R���"���  |Q_�`5�5^��/�/3Ѕ�����'l��K�ݰ!�|6\����T��x�}ffB�)�
*:�=���Й�h��UoVTVXeU���;�C��n�3��&���GH����v��>�+�!I`���W_釗��7���Al�RR\*�^o�2��}.,,p~mo���(qE�j�ܩ�(ոyP�M�4�n�ͯ<�O���ǭ��]��`6��6��rږ6r��k+�v�Yg9��X� &F�0��Cf5�@È*.�g�G�.]�=��Mu����팙��4�/��.S�N�3������m����7���"�=�"�;f?t� A����7ߜ�F䣏>�r�x��K���\�t^��b��dqq�o�A�h�2kj��5�]�d���a.��ݶZ�evN�����q�~�=�����Z��6p��nu��uK�$I������/k�:����2�l͊�v����>ceC�۬����e�"U]nPҖ�� ��d|����^�X�Q��C0��l'�=������Ox�K.=}�fl2��K�?�M�����q�V�/�~>�{�Y�4yK+,(��+����a�����+<(�t���.-�S�C�h�|����S3f����ټ�sݯ����+�0Wªƪ+�پ��yG����"pܱ�)�NH��8�)r�I���3��'|�T=�ӛN����Ay��a����� �.��";��c}Բ�^
 ~�������M�:�,�h#��]�P�I��P���s�x����E	`�`P�@�m}]���)�9�݂���[���?��~�1f���3Hl(ҸC����b�H�T���֒Q��R,�]Y��Uu{^�w�q��u���s�1�(��x��7�!�@�,=����_����}#�t� �E�:0����
k��T7쨕��Uz|Y��fW��l�Q؂ x��O?/F.4y�Gl�[oXY� ����*�?De�ߔ#(MaƄg,�OS�5o�l�v�FlYק~��ޖ0�(7�'&0��5j��!���Q߳{�,G�D�x�^�/� 
��}"�l�2�xR�|C(��(�h�7�͘A�mq����8��(ВQ��`��H��.�mvc��Ӓ��E���A��}/HI�?�A,��G�D��"�6��F<'p�;l[�Wa<A����C~a ;�5�q���(v��%����M��I
�_�[co��rT;���@b-2�1Cy�%�O~|�������SN�����z\��z�DfJA�5z�굒Ãl������e�����ɑ�"�p�_���Ԅ�(���x�=[���VT6��(���x��F�h�*�PO����ړn���>�;�-�%�brj��t�7��k��n����������>ɦl1��J[bM�p�<�6��A��v啗+\m���Mv�� �U�ά1���P�Ŷ�ldD�a�)^����@Lp��=�1�;lk�����瞷�O�����[����q��HN8`� m��>Ӆ��aB��+��t��d��j�e�vm8����ZZ8��
r¬!�K0�aj��W��c���}.O<�d�%u�+&g�H�����Y��r��v����R�=��C6v�X�sϽl���*��(� ����C8Mm�-[�Lx'���r��|�=�u�ό�Pd+V.���L�񏮱�����N���Q����*U��ꏘ=íي�dP&3+[�����L��T�[�ҩg�"��K�[nV�u��s�2��1�U�%}eH?�_��w_~��M]��1���>�~x���_u�O�v��f{�M��7m��|1{ΰ��~�Ru�~饗�p���+��^�Jt��A���5B2-������p7@I�S*b:(Utv�E%�:Ӛի�($�����l�]wr��I�'y�����o+��&�ܕ{F<ɓ��`A�pÆ�	����@���1���	�"�G�:�i[M�����;�
\:q:$h���#Ghjjm�d�\Wh���Ӏ��6Wƃ���>c�B���uԝ���>�y�u��Hx��t0D|�,���q��G'P��S�/��D��K����&��I��Q����I:<�7����_h�tW�z�<cT,�7�eH3f
���F���M��NŃQJ���(�2��p�����)�*g�<̕��A,/Jx���Y~^N��������D�3�P7�ަ�$�Ȱ�Am�Y���e���Me'�g�@�p>N��ys�R$��2���
�7@����?I�����s�K�2X�_��������7�����[�JPXQ�0��_z��'�ƤJ@����8�	 xFl1N�DZ�G%=�5���=��v��3����H9#��#;�e�H��oI�o"PǍ�O�e�>��)O��qS�������c0���/��~�ӟ۫��n�}��+.�H y2X�!�L#�L�Ca� 9�"�"�����;� �;�Na�%��l�	4cЅ6���%��"�y��x��[jK�` 9�`��H�o</�1�|���w|��u��g��]r���և�o_yՕv��*Uf�2���p�d��^�{��ڵ���~��좋.�RTX�8�=e��v� �=�}��6�l^H�P;�j�����:���.{ꩧeĝ������޾���]����뼞�	��Mn��v߄��7��3J�>��o���	MZT�,���vĈQ֯t@��M�{7tuɐTY3��YcS��];}��[��w�X��O�Yf1�0X{�x!�cV�����=�塇�h8�@{���ݻ�o�'��YF6ab6��>�Ï8�����9-_x����.�E�ڸq�Y]C���ٕ�]iGq��xOy�(�'�8�QY��?I�����J�2���-�?����O���z��Oo���Z7f��-��J[�t�x=�3<���[�)ʘ������Ҏ��ۧ�oh 1��|]�+���3fl2��K�?�M�����9�?��5�<��i˗/�]�v�*�Q&kP h��1��Ҁ}�GmvN�"9+��w�\�t���⍝��ΐ�s��KS���!�YT\W_��2]�H�m��V��_�lӧNw���%;�o�3k�o�w;�' ��C�#ߘ��GH�=c&��B�{�ˋ���་}��W���7'�>�� 3�JGC�QJ188<��),L�� ��\hRT�v��}�
�0�BIIkm�r�}F 1��EQ&y�NO��!iǴPB�Q���ka8C�gt~�C~Q!��O�7P����)y�2�K��Un�F�1����Ѭ��~$��੽�[xO4�wU�*[uc��������!�gK�	#��m����"�pEM}��7|�(�2b�ͼ\��
�L}�3W��M�愪���.=����}6Qegfz��i��JQ�S.�_y�*��b�f̟�!?p���~Ř�瘽�?>��c�����qH��{~�ߐ�	<b]�WW{�U3P�<`�3�q����a�3��J�1��$=�w�mrO�1o����uA�|�h �����7�D�l��K���H~G�{���@c�^�7���>#��R$���ݒy�L�h���{f�|��*����|�6�,���F3H�=�l���_�ǟ|b�z�+�;��[!md�����^�uت�<��/x���z���|OY���}�E0�Ծdh�Y،%�e� �S������G4c��'!Gm?C�U�	ϐ�&y�]Gg��}�w�{�\`�w��r�ol��1�P\R����.�'N��Ԑ���/|�U��&=f�0�~(����b�^z��x��(�h���x��ަ��@JO��+ �U�hv.���ۢŋ��SO����w���I'��4R}���7\��{ 6�8��s}���"�!v�c�8d7ۤ�u?�J���w���4����.((��e�z���m������l.յ�bf	�h�oq�~ˀ8�����6�,���A�ީ�ef��>�l��/):��.v��b��e��/��a����g$�H��1��X[]!^�ɾ}�I e���q̉��S��f#[����v�E��A�*Y��ڃ�A�hMQREk��_��1�����z��'֟Z�����k�$�N>�d{�ٿ�A�d��u���5>���ӏ�L����`�/�ZO�'���S������h q>�
�ǠI�1���Ͽ��]v�e���	��i��@�+�?��G����@�ǰa4�N(

�1W-����>ÅE����)���s�M爀$=�)���~���!���;� Q@���|�1G�h��u��@��v��ҥd�1s�y��2��}W:�(�p_:ሻJ����_����O�O�¨��Śd|��>�1�N��{�ܹ��L��Ά��8�JYIN3= t��K-ڠ���0*���"��� ������.W0Q��X���6C���Q� ��L��##�} �E�c�i{��c��#: (�=�1�(_���{��Uy�6�	���
/�4!!�(bj�ޣ:_1��Bo���iom�2��H�-�1�Qq���,��=��9��e4�N}���s�Ï��ʸ-�Q�|��<1j�i �N�A�)f�D���mhAI��٢�p�~��N;UP�ʚ}��E騴�Hg� o҂���xq�F�ʠ�ށ�}�Q�H�z�\����R�3�t�3�Ƀ+F�D��WF�Z
�6��5I�IK��
�.<>�˴�P�.�t�Ŏ2x�G>|�P�}�A"�2G��&B��D -����|��	�=��Ғ�Q�1�08i# �[���fA���Ka���c�:aW1�,Iƍ��Mx{���������s��o~�~��[m�9~�pUe�m���2�?�8Qn���Q��	v�5D*K�� ��2�0f��~
���7�HRZI�����p��XN��(kdb=��/(�ק2�4�����AcҢ�Kշ��~����^���;��h��Q�M�v��G�e�^%�)�����r;�{���)��d76��[�����,�397��s;���?��.��R������v������ 
?����ښ��l��*	�k��5T�c�̱�;���v��_�2~�����o�������F+�骫�� �!�����y�Y�[n���~�m�񠟡>���u�\~��f��'�x3ᔧ6Vg_�����R�d��l�n��omV�9r��z�-��i��岌:g&��]�A��T�n�O�D���N;E�����~�;�}�{��_xP}����V�Z#�ɥ: �g3_{���f���om�}�q~��nV~'���<nC��� �����^cӷ����R�[-[m�85�2���x"����[������hhW�h��n�W=����g�|�z���>xp�wYAQ��z�������[o���>���>���c �+�u>�Y�����s��ީ���&�����	�?���ւ9s���6֧�%B�w:-�r�A9D1ǟ{��9.��{�=���/\�3"���]+�RAZt��I*��H�8��뮻�~������������.�gxo"����fg8�b���]���aD�k��%��'����K�.��B˗-���*[���V,_m˗����\׮�е�j�����e�h���X�l�uM�DD��F��i��+V��/�ڢ���I7[���Zm���ưn�:u�k�7�Z/f��ͅ��P8P�xN�`X%*�t�К��0�n�"n2���Y,��afF��RH�@f��#_�]�q؂Zy�kZ ,���-�26��X�Y�7
�0؞���p^�`Gf���.Z����]hO<��]r�ev�I��	ǝh�}�8;�ȣ��#���<�א�<�����|�M�9҇��@<��g���U]Ya��\��_��?ng��=w=�Cm�=��]Ķ���+k׭��+��R��(��9����/�w�`�`DFc��hOԃׅPBlӱ^y�{�3��u��6�Ŷĕ��2Љo�]�=p`�M������6y���~ʌ�g��\w�|�%K��+ 2".!ݐ/����@�D >e�؀��D�ن�t���Q����w��uCpx��� 3�$.\~ӎb��'�1�m�40F��gĉ�,B�71��|�8�;�a��5H�Tң�9�h��aNG�1�A6�&)nW�p�"s�-	�b�(˒%K%�V�[��.Y�v�� ��v��նh�2[�l�Ϣ���r�k\ɓr�M1�\�O�+қ�<����x�����o���G��n��N+:"�3�m��@`ժ�n�s��I'��u�QB��+�|�+@{��`���%2�����R�ڲ�+�?�i�ʻ�r>���}�4f1�%���1iP&fu��m1��G�s��{y1�8+���� i���H��+.��ȸ��Yg�����#MfY�D?�YQ���12v�v�J�������d����^�މí\b�:fԠq��>� n������+�uE�E^o�ǚX܄Q�,�� ��f�@gXۚ��aU�f�<z�q�=��{�\[Y��ZE�Z�j}M����Z���E����]�^�{hɇ�B�b��V߾��#@�[�9�)����e 'h�������?�y������(�&���&�k��m9�,rԨR�D�!"�	��MC�e7#��L@�X��;ԨL�}:���+ ���M��w�߷#;�x�O< ��@m���B8��O`7�;`�q��	C)����$���/ťP�Q���
w\=
թ�K�f=H�ee�y��Z^>kCB���B��"��W��ߤ���7�)�{ȗ�_P�
��@B^����
��\���Ġ��-|��(��gS�i),(��;=˲��p�T��������
.~��%�sN�!�RÚ*����M�����	fup�`�taQ��Ş~���9�5=[�	Ǭ<�$�$��-;?\eT��S/��AVY*>�q�ڈ�tws\�|��,..}�������駟r�&�.((q <Fgo�ô��;�9m�g$��Pp]y��g]1c�1��,J쩧�j_t�+���[��aC���aL�Wl��n]���5�N�H�'t��D��ۨp 7�kTp�x�w�y4"�����wQ�,Ƌ4ҥ.Q��BaEQ劢�҉���~���B�� Q�����~�31$x@+�@�7�$qb}Ő�N(K_�@:���M�+��Dڠ`")m�t�c�y1B������X��C���A��kyF�w���ʜ�!^0Q�7�|�}�=��U��f�-ϟ]{͏�׿����3�~p�_�e֘`�R���jk�lQ�����E3��vu�I���ĉuͷ�˖zy��r��[A5H,/���@a�����S;�����o�~�\7P0�|���������W�}�����oW�Y��z[\�¦�PD�#h�Ҍq�Z���0��~p�evҷNQ[��ۀ�d��u{�]wݵv����IJ�c`�4 ʄ!/fo�]����n?��Ͻ�c��?��C���9��ASn��H�!���O����׿���[ߝ��]!y�7ƾ��k��{��s�mv�?�3��/@_;`=��B{�������͏���a'ý��Ǯ��j�_/Z��3�[t�&o��ul 2t��3>���v�]w�P�N�2��`$��E�X65xO/K���+�52*?mXcW����U���fi�]�b�{�ݷ�%�)�맟}�>��C[<w�5��������������y�j[�&#55�E���s��t/��'����@/_"����E�Z��Ѡkpo�B�o\�o��%�q�&�Z@wWw�!+V](��Wo����b@���P<F��Z���&����N�A͕M����3�������������٧�yG��  ��\X�NB��+^�s��p�m�������ac��ȹ��<�cp���{��*���T5�V�b��ꠥ�'�1��a}�H�@Z))��+])8�Ă�Ƶ����MhB]��p��[�8��BG�i�Q��,O���=k�R���ߤ�^�4�/�D����oz�w�7��ȏ��1�[������f)�R�8���ЩÛl<�BC'y�<8+�]�H��ןa2e���---��C��0(�����>v�&�wP����PxɃx� �ɕ�(wl���3��_�=���V$�w�!n앖���G�)��w���I���~t�O|f6��f$������f����;���0;�yG)̠U��aKS���we�:[�l��R[�h���+�����P�<O�E����u�{��>P�pG|睷�`�+V��P�p`���(xą�|�yL3�M��D�7�)�6��# ��?�e�2����/��{���{��<�\k��+�p�[�> 3�ĥ��"�`��1C|�"�׆�z�Ff޼��ɧ�Z����d<��cN��ٜ�g���!�1C�9B��K�w����r˯}㢋.�/��8��[o����^���?�k�˟�λn���3��v�oo�?��n���?�w�&�Y�M�N�"Oy����^�P����\Џ6M[jkmv�|���~a����v��TI9�wF��36�c���%����	x*�W��t'�Ao�- ]��6W�uםŏ�ʶ�f��V�����e��w0v�d��7�;����@��?�AX��������E�6M�0�t�	'����3)��pȋ�o #v����窱^�u���v��h6YHI���e�/��(�a�Z���:����=��� �����A�U�V��nO<�]~�����gdn��0[���ؽ���9� 2��v�e{wo����Q���� o�J>�)P{w������m�V��mE�#Kmlͪe6�<[�r~6�}2g�}��6��ϭ�����d�I��Km����+��N����oq�o��g�=��@|����k �HK�E]0��xe��������ڵ���jk��\)��R�%�$Ku���Ih�>����ᏰG��]����	l�����!���#�4dW��zD���b��f7ذ�A!D�YCJ@"�b��+���w��o�ￃ�#���5�2�7� �F2xZ����^��h�	M��TJ��f��ÏdM�.ݸд����w4[k���$=K�w��5���uעM��w�y��%_ʯ�[�@�VRum]��&��D'����u+�UxQ'�A�^Ɩ���!�]t��a'&�PP����w����M�Mu������=�]e�Qح�ݝ�pU/�����d�̐��wg*�q ;ܥ)Ї�K!�>l<�Q��hnM»-9�zR��v�:�k�H��.�Sa�%�gYc{�5)�V��$�)z��)~TH�����NVwGw��+㪝�[Eo\=Dk��V\��Uʭ��.G�a܋p[�Á�B�g�<�3��1Ŭ	���O�C;��8�;M��G����{�R-�����`��e����/��_X���6v�fVP�cS��`�}�t��_~o�<����W��±�6D�X��lW	��w��v�߱�v��v�m7�޹�ؑGiEyVX��:b��^e	剰�����>t���p���|��(�!P�*+�dU�!�x�Rw	]�l���/]�D�@��ʻ���]���ŗ�W��:�3ŷ��%����5�=JnTvb�b�4�eJ�F[f� ��U.�� 	�p9B��m��[{�G4��I��>�1�5�(�`̔��O�yz����ϻ��H��|?|X�%�S2Y���E�1�S.����~fO��l��v˯i���WRt�e$�Xmu��v�e�=.�e�����fZ��o�t�]s�v��g�ȑC�޳��Wyu��&��x���u���>��~v���~��c{�m��v6]�>l�P�6}���k{e�`�������o����0��Y:�l�D=��a�L����'��Vt���`���RZ="!�IU����z�3$|�?d����"f<���`�n{��,�3��@���v���k|�3�nMM��/߷C�0H�Ȁ�RkV}�̤2����!GCT�TZ�dv�d3a��96�l��dȠ�oS�L�����՚M;0 �U4�"�c$m.B�b�ʲv�r��!c'�L
tu���E���������"���
�"�9r��Vdcǌu7�)�O��7W�H�xH���,u7�f\q��8�p�I�ջ�#0y�П3��DS�W�Û.)S���++�--��f�H<�x�}��(�*���3Ǟx�U{�\+Pj[N�b[O�j�N���
�[C]�͟�����틆�a�mלrТ�[:��9\i#�`������O_�г�ɑ����D��wC�7��,�a�F�q�ɒ��9�6���Z�&�Z���3�/]���?����n��zG�JB�8!�5zuo�8K��@P�P}���������L�?<��FŨ���;�(|pM���>!~4�\�y�J,!��~��o(`�'�@^�̔��٠�%Y4KN�P`G#�W��3*�L8��]��4�$��Q��m�SG��*!�� �#�10Rs��E�iTGZߚd�2Z�e0$gY��&ɿv�I�֩�m�F:z�hu�ɠI�����FJDO���%[Ss�:m�J��5�Z����kT��f���]�[�{����N42#�ɧw2x�A�[u�!�]Wr���8i:��u���E�J�E�u�xF�v�3
�κ+����d(���.6l,cSe�>};;�m����!��]�$�+N��'�T`�i�8�d�)_u$µMg��ݡα��C8��m�zMn�c �N'32����Ε^����:ߢ���Y����{I��K
S?k��:{�,w!e;���[�f�����2z������^���/H�h�q�︴�n;�.��`�����lkh��-�7O�u�.R(~,�F��W��x������ݺn��F��7���n����r�駺B����L9�M�߉!�}�3H��I�6�h����Z�y�b�14F���kiR�O�h��q�%��~�	9ԇ��A�I3*���;4%wE#��+�(�PD��dv��+奞iܤ�;~�B܌ ��o&d*ϣ�,e�`��6d�_�� T�d[��t�}�멄 ��d�i�1��ѭ������N9��e�|�/n����.������ϳo�p���O����cF�_Jl�=v�3v�>���;�=�<� ?~��u�����8@�/\��f�|�f�=�~�aߊ����]ʓs�.��"w����W��~�{w��|�b�r���U�yb�@~V��n�wX�1:�	|\VV��-��d���q ���tӍNʈ�"��邏N��:��:���lĈ��>;���z)�2�A\�]���=�½l=(.3+@�?�9��6i�D��eC��2<Ə�$�h�x����]=j������#�=ކ�m`!~��z��;�������a@�O.�YT�12�U�2	�[�[Z$Q�e���J�,a�k����勋c���-;̔�,�ܬ��48ߐ]E!��44Y?" �^�����n����^S��mٮ%�lTv�U������l�䩶�����[N��2���s_;��í� ?����ڐ�<�6�MJ�Q̸���a�a�Ox�	�(˿zO�������ob���3̀R�I��M��	�a|@J^�:�4܀�L�#|������
R0�G����Ď� �F!6d�F|���IޱU-]T��X������:�Z1GIE�e�4��.����������6����gA���e����a�����b2N��P�e�H�o�үߝIY2l�2�3%CQӭǃ~�����ѻ����6�L�n�c���X�4�R��-�|��k�#�ڄ�ٰ��[Z�PH٢Q�5�gZ]3�[�57�XkK��W�2�Zd�t�ZOj?y� #�Y8�*t($'KI&E�']�c܈�d� ꒑�ڑ"cH�Iε���\�[�����֥kgc��+�5��iʱ��\���雮kn�R}gː*���!���.��;�к������%M�\Cu���vڷ�k��%�#�Y h��^/J���+�8KA�h�#��I	m���'ۤ�';O�C�2��~���h�+���Gގ<�Au�1B/c��ㆃ���Kl]�*�C��P��3���\RR*��&Ցg���Će�E��K,�n�o� �����w���V\z0�N�~p�'�~��c?4�3_�<�Hww��C/�'��i��g�$� �>1.t!�7�gv�{�-82,Q6�h�+�%k[ȟ�}&%{=>�0� )�A̗�����ϩ��4J&q�"���(�|�`�G��<��#-�!�=G�P�b� 20�LF�Ɔ�p�3�59}�a�"}�04��%҃M�+�fr�^�{�7e���g�a�����R�|�{�@cv[�d����	u��K/�A��#�8����
��o���~x��G���z�!��og�S�p�>��^ַ�HSʉ[���-�'��R�*1�>�-�U[�p�V�X�O�E��_�]
)'#�3���Nl�|�Av�G�әg�i�\r��A�����_�]!��c �<� �c\c��^�y�@aWb5j�]|��~��\`�]z����:�,�:���<��"������;���g?S{�M�lu�u��F^�Ft����8l��L���!ʹ<�)|��ﱇhs�p@X�uȡ����o�v�QG�Qy�1��q���<��|#�8�� ������ߢn߸�B��|�0��6+=�j+�}K��kX[e�����;�f�ﲻdc�(��/�6ґ,��Ͷ��6[��ql`n���n[�n��X�\���/R,��H� ��,�����N��
k��V�L�o��"�d }�@�+9##3e@��3;�X�:����_�%d6��\�%��p�7���EAwOK�`ӡ�w��w/�0�@�B#��I���1�g�����<�
S&��e��.��M�R��zdHd�萡d2 ,ǚ�2dXrZ?	�J�L�*QG�/�0O��LK�hC'ΰI�`c��aEçXN�X+>�n���jw:a[+=���m���[Ѱ�-��hK-n��Yր1�;h�ԻI;d;r��x��6i�m�v{�$�b}Ӟ�O[���2�JU�bQ��RuM�)�̤B�N���g)�������Ι2�d�� ��.R(�a3�R
GYWj���"k��o�V��e��Yj2ʺ3)��2K,{�D�7n+5�
d���n��Y��)6`�T2q++�|�iM�g_�i�IyVP8H� E����U�(���3���ם��2R;1X��ÅT��&��!�����N�-�"J�{\t�b}�?�SW2\9
���OG���s�u�Iiƕevذ��A��Y�lt�'|����O���nC����n{�wm��
klhN9~R>�1��R�[�&�$�����;��}��(m�m�?��Wb���a݅��F�
WT�2��<1�.�l!0*�r����;����	��3�/��F[��<p&�k�B��Q}0s��p���P]�e��G���S����'8p��f���hd�s�Op�w���`SʊqD��\9�	 ��|��]Ǆ�ϼ��H���"����(�����q�ܾ[��z�;���S�,�W_}��x���a��+���g=���z�PF�}v�?����w�cV���Ǝg�l��>Rr��|��U���Yfț�Aȟ�*��f�h�d&�+��S����&1q=��@�pt�w�/�0�o��3[/����K�,1²�*���ZG��Еg��s��@�1(�}u����"�D�]�w�M6%�������Ae6n��b������Q�٘��l��w��7��#Ҏ��A��7�Ct� K���ov ��3�� ڃ#��U�U�c�2�1�0z0(ٶ�Ck9�h뭷��'18Y�,Fܞ{�)�n�%����9A�;�p;d������	�&fr1��mт�����|��}�M[2{�u5�[��J[0{�U�[k�jG��V��s�ټ�󬩭�v�}7�8n�U�Xns?��^y�y[�x��p�n�-�����������Z�,F}����G�J����k^�M�}f|-@B(Y�5�]xhX(1�!G8�u?��L�f�%5Y�A�;K�
B�@��=��tl��9�e���g� ��()��a���	�΄��%A���%	��>�/˅�wb<B�� p���}��QB/����{�5�nnW�Sd��-)�������Q�R2̺�K�S�zkM�B���fYKu����[W=!�z��7d*��I�o���6{q���i�)�=�֓9�:3˭95�VI�^Z�f52������2&M���o��m��!��G�6�aS��(��Fm���������O�12vK��l�:�2�7�q5�ں���%G^��7eK�ȴ�k��ҧ��$~�*���Q�F���-�d���5v������t�>���;s�֖3n[K����j)#���ͦZ�p�%��d�6`�)3�����֖?f�ec��GYΐ�6HFR�����'���z�V�k�Ԥ"��Y��wf[KG��l7F�L��̵�Ѻ�٫��u��)u-I�ڋoڧ�[��%��s( �|y�ݱt�|����9�lJ3(��z��dd���ZY��,�A�O���Bc��:�ceE�}��B��Oۼ�K��o!c���/��
��O� J6�Oܭ\PQ���}ǅ�ę7o�o=�;6I��(Q(��	���m9/{�s ��W\ɐ����(�(�l+�25a�?��-vBc�oF��1A�ŀ@�G>H��@��#% ��d e�e�+V�'�S�c@�P�A(�����F0�D̗�h��F���m�مc��#��W_����]"�('�I��ph(u�s��G2�Y�J�E�B��&�N��g(���8c�&nȄp�R�����)슆��䏱�����7��@qfC�O>��������n��n��1V6`��J΍�����و��sgmM�U�������W(7��R��IR�_ ϻ� p��1<0<
�d��f�gf����SN9��G��3��cƌ��$e�H���$�`=t�Ω�D�x^��w�T�������t�����EE^��k�`�<[�d���PYU��X.Cn���R7�0`_~�eoӫW��r�# �(��pg�F��x/�%�1p����ܐ�9s��t����/!�^��d�F��[o��e	m������ض���^F �rlC_����7X�h{��h�z���z��:�5g�}���x�"�je��^}�M{���w޶W^�^|�E���gV��²�3-�w}�T�X��� o���s��#�Mh_�61޿H���M�K��dT���7�6H_3P�������S���(!��)�(:�#�I�$t
4ʨ��(�t��F�"XYk;���<>�m��FEx�s�p��(t�_���"��|�x�t%*9�]|�7\��=�=卝�w4���z���GG�=J�NON�9��M�ֆM�n���h�e��4�J���jG+����i)����%P�YRAK),����֓�o5��sq:[m줱6l�p��o��k�l��z[���VI�^��cqu�ղaAQ�%��N)���V���N��b�:{j����o�����g��d�*k�ȳ��[�0&�6�d)Ń�2���9]���� ���
�=��:2�Ywf+1نL���o���*�M�fecFY��a�]>�F���&ﹿ�����<ՆJq0eK+M�N��O�aC��ڎT���ޖշ������VT7�\m����VֶۧVٲ��lJ���D7��-ǚR�{��ҚiM-�Ԝ.�KU��Y)�,C)�p����4�%��;��
Yv�@kk��È�����*���|�KP|y�yKm����3#�J|�{��Y1�m(�)�ʐ������Yw0��e�V�{�}h�������oР��W����ȑc��C��?�Pv�g���'({���y�=�1�2�R��o�"E����6�>ʴ�
 π�{��]I'���]��G#`��T�O����-��)GW����\ ��Y0<P���x`�!�6�8#�x����X��Ha�&������$}OھP[�2�?�J���.��z]y�3Fӡ;�1�'\ˠ;�·�_�{�јv��5��(ǐQ�%N|���̼CcA{�a1S@�QVO�2�wPc��]��!�}��O�B|�f(�؅��+��ٿ�@���R-�⩔:d�m9uK�5�G6D(*.�f��zź����Gܰ9��D�9F=�(��55������)�	��5j�y\lW�.���bD�6���~�2�v~O^x>0��n�xn��aS����H��#e�<�&O�d�&Mp�m��1�u���k�X����l3�Ҏ�����U�ZC�h�{�$�����:���r"?X�Ħ��Bël�Ρ�h�`Ƕ�n�|��S����<�e�]|Fz��{�A8�Ol-_+��ȵ�]v��g��+��"��N��#�2�K$�$+Ey�ij�z��-��d��K�����X�Y���X�[��@t��T�y��oi�*c�w�`�Ǩ �w����6��b|�<b>��GH��
�\c�&x��/�'Ҍ��f�U}�n��=|y8a�?5��U�VM~������R����*UdS���(jia��P�$Ԛ��j�0jUE�h�����"��=���I�h̄>���/���CK��h�#��o����ܹ�GS�=ֿ��
'����|Pn�/
��>�"��|��=�!���ş�x|�>�i�x|�i�c�Sm�]v�ܼ����l��
+>�J������1l���]�O��m�]���v��&찭m��ζ��;�ح��I3����m�3l�6[��-7����X�:ҝ��Ɏ=aG��-���F+.j����5n�U�_�N>+/�r
�,W��BU2\[D�t)��2�RTGy%������+PfE�鈊,� �rK������<ɆO�܆)����:ȉ3v����a#�L�Ԓ��=`��J���ʐ!&z�:%��6h�p.CiĈ�֯d���%ggZ�p�Q���R�����y����Kga)[�sN�ޜ�|4`����0z�ujI���kez���c]�ٖUTn��C�p�h�(˕!Q�kɈ�V�gY�X�q6}�=E۝�d3)��X٠r��~�]w�%�g[�λ�l���hu���`�X�t�=��㮔aT����Sr�Z�-���ͳ���R���]�������vY=��TW�Ȩk�B�+ŧ��imk�r�6~�X�lڴ)���Ռ��=�����Y�%v���:Z�j��ˑ&�PdY[q�QG��[^>H��07~�+4�e܇P&ߞ�����l�v�5��p��;�/�xO�`���<�pqcI�嫱��Fa}M��)��,VU�$Y_�6��%�M�<M��^�͎@a}$8B�h���d)��2�Q�P�e@�0(#����,+;�뎧��2��s6@�uL��6\IS�gPN8���H��%�=H
��P�æ4���讇�;���@��J�U��ya���  ��l �h�������'u��3[�E~A���̞�Y��N;ݶ�z[�Ap��1b�xd�oC?�"�v����e�u��yp"]fl|-��/�\�l).P{	�Q?�"�ls�8Fy�1�q�_���
�R�U���M�>�2��4���q�~{�ԁ��q�
����@��#�:�~��J|��36�����d1۟S�W+$�9�99�Y�&@yv���8�︱�	�X����;L�媍�a1B��~FT�d@^~�����=�WT�����z�!~�Η�-��Ζ�{p�Cv��.t7���f_눋܌vvz�
���O��9�}�cOk��l�m��N<эH��l���F�pv�e��,�c�VH/�l������'��z�A6V}���c�=������	gge�a�[l���j��V��80��{��7�jhU;L�eHF�H���2���T�\ks�M�J��� �/��a�O�ͫ���9s���[�O�bs?���:ۺ��߲�ޝ���q�xuy$#*�<�J��.�K<ҍ�#z���b~@�{�o�&|>̚��n�#��d�R�O�~��b|��˵�_b��`Y��6����eq�W(y�B�K�\�n���.]z�m���y��p�)*�E��樃�E�N#I}��"�O'L���8_6�\���֗QL����A�s.j�E����x�?o�l?���3��h�|?�����o~K8֪��FR{G��n1RG�t��փ Ρ�)��F���xtFt�((�5ո���(��<ݍ����%Ur�]¶���?�H;�g�Q���Oۣ/}h%6�����W:�rJ�Y�:���V��-��o䐗�a�KE)5�-��N.C����[�Q���n�׶�{s��&y6�,�*W�Z]��Zh������U����G��ft]���}S3��Д�uW�luv(���K螖�f��ٮh�HI���R��Z���s
n�L��Ҭ_q�5�v��/ڲe�e`��Rk����:�_TbU�=���Fu�j��*_{�շ+�lܠr,��g�&Z�u���VY��I*�2��H�<ѨPFSv&M4ي�K�������E��.��+E�P
�P�p��U�L�|SS�`������h�5k��z����a����i+�|��
0g�,�g��}7������f�1G�.K�G�p:�?�D�؋N�]v*�ڙ�=�n��z�	t�������	g�L�8QFz���q�/J��aå\��vg��'��W^�QcF�ĉc�.p�S3	�y��7��@yB�ekP�QI����J����֮�uA����
O <��}/��x����m�����&�`JP�Q�����[�+��S6�`��t�`D�no�!$�FYB��&/F�Q�Q���d��i�1N�y��3f����x�MɁ���)C,[PJ�|w��O(��A��55VUQi�j�-m}���{����)��{j�[�a$C���Ě�u*[5�YJ�\I�g�D���v)߫܈��/R��[x�wq	dGɠp�k�jw���qC�;����Pn���?�"�72��!���^v�2(�d�D3�f�++W�[o�-Ȕ���&��>�qM�[/K#}�U�*�Y�k[�-X4OJ�*/�^{��.��_v��6L�j+{�'}6m��H'���K�V[M����%bs ������8R�6�b��s�4��?�v�pa,�q��e�0c'Ht�c�v���K���������:)c硇m�x�kd\r��{�/�c��ʰ���<��I��g ^����>�o{�~}˯�8"�\���<�T��/~��<������}O����+���.��
���%O>��xc�Sğ���d�na'�r�e��A�_��3 �ƁO"�  ��IDATF\b�}�׳�>���ٳĿ�v����<�㶷vٵ�^g���#��n�?�n��&�G������?����w�/��Q�L���0���gu%[���WJoI��AC�g_|�����5�چ����w޲{��>���ˠ���~��YS]�]s�uv��n��=�A�x��c�rJ��C� g �%2����ϸx�l��b�O_	�����aR��������N���[n9��x|��KASsc�ʕ+����T�b��	�7�(\��)b�d5�d1n��=Q�D;E�6Uq8,˟z�Ҩ����;���Ҋ��^��[i�Mb�B�� ���N��ib���.Fv�Zu�J�|��x�X�Gǟ+�J�KW�=Iem�:��'+���'ݧ)��PK��(���z��E���-HQ���Z)i���-Q'�%᳋�����K�/0����(�X�o:k�8���%\��q��3��
��o�.p�̅ၑ턗�pOæse�zx��Qdex�8�{�=��ӼG$eq�����x.r�lА��PN�8�	�	6���8��Q@Q�8�%�m��A("�RS�]��[�-�a�\��ab;oߌ��Q��$;�#��m�J�g�nO�.�{�X+.mM��V��f5͍>֯lPP�VWy��龆#I8�#�ū[�9z�7��-���f/ݨt)�2P�� ��,	J�Z��-ǳT���F��e f�3^�:č2C�`��-j�d�;%)��d��X�B+��3g��a���}�Xuly��"�Z��_a���)6vb?[���*��IU����`m��uv�SZ-�Rre�`X'���D�Lu��+uN��e�.���,ԩv�`�%Y�:���f�7BJҠ��K�"�L�|�թN*�j\!��4��n{��)9�*U�t+P_�?�ǆ�I����g��:Z�I!��;It�����9R���Q��m&S�q�RO��P�釟ᛁ�o��-���u��m��w�b5�>��c,�y��Ӥ���� K@���bN�g&�WL���ff͙-�p�͚��2Q�ؓ)p���I���30�����$�af���0_|�d���S9[���P
Q���A�B{�
o���6��1Wh�Ւ��Ql��ۼ�F�`4���[�����>��l���WUV[S��N�)7�'p�m�A�m��_�	SȐ(�Pr1���3e�� �l���2���*d�2RY�g8�vm�d�~���������y�F��U{�=��d�8�BT+c�G�;�(�L��dQq��H�Y_̵�v'�u<�'��D��,<�0h��d��իW��O��vy�cb�]v��.����£�KeFi��w�C=��r��FΑ'x�z��[��{q��z�؆v��edE�m~-�ܩVY��������>P[	�B2�pǄ�hC����s}��#w �@bV��ʪ��< �	�R��&1s��7(��<���{������ܨa6��.�믿Nq���l��*�g�m��/�r[m�͆�#}�Ǝ�%�Xw����zͷ�g&7��p��d��
ۧ %�:a����6�xk�>аx�"[���;���ݤ8�@z���sϵ��U��F����_�����S�c�>��M�6�
�rշ�Q�Yl����=E�����k���C��^��s���v1|�e�t�H����l�n�Ѯ��U��f>b������:��/^����?x�w�<�['Y��~VQ]i��Q��⥋7�3��:��߳Y���fC�[���6i�D�_f�_~�u�m�=��㎱'�|��p�]6{�ږ�$g~�����
���ծ��'��[6n ,3@6�$x���;6�G~���3�O!d#������/�'$?7M��<�b��~�������d�R�ȭ�����O?���ӷ��	l��=l��=����kkj����J$�7���Ow�p/��K!M�"�Y5/�MR� n<��06��lJ�(��IR�{�{Ϣ�	ОήΤ��F$�G|C�og>	�1]��?	CJ�y:��A��8 B�4�L��q1�`p���r�~�q'�KR<�F�z\���$�>s#Ii�r����ݙ,:ykBɏi�6�YO��9��2���R�o��-���M).)v?jAuU�w�4�ի�xG���<�[ZQHD�E;]J>�pKA�WV��W1�C���t����pE���.9�֭����[��{�a�������%����|F��k=�e|�	������Os�o���v�~�J0H�#'�3�D��G=2ԆI�>��Sv�wX��I8v����c�v�u�gK[�l���/�jO=��4c�]}��V0����ؓ����Xv�1�Q<Җ�ĕ���{T���|8���Zա�t�7#d$�Uw-�'���VѮJ�et]�C;s�"IB�C\Uaҝ��p�Oʳ,�?(5���62M��F_+����xA��s*����t�y~IRf� �X񤰣�3r���n�~R��a�J	-����[f^�-Y�Ԫk�']��7Yy����"�;%�V��$��]r�V囤�����H��]+UN	�d���.|h�R�12�zvieI�g�P'�4/����b4y����&#�=M���ly9�6������Z#���oY]M���c,.�?��;� w�(v#�lɲRx���{ۆ礠��ϴex�J�E��Y](�9�y�k���+�~���ZF�7^�
�[�`o�|�^��1󭙶�:|x�Uty�ɧ��?���&eb�}��}�g�0F�����W5}��V*���DI���#��G�D���>�I��8�XV����%�����kyP ��dk�X_E2�{*��0�A��r�v2�|SK�2r���g�K��߿��T��G������:��&O+#=Ǎ��2rޕ1 =]�a H��zHG	%'3���k��ؤI�mР2əj�F�@鯪�1'Cb0@'�D)��->c�b���}��3�����������ҍ�W>�\��c��k�]�΁���OAQBl�٭��>�о}�I���\'C�I���FЁx��X��@� ���~_�����:|�P�R2vu��Hm �3~�+��p/��w޹2vX�p ��/��q�]��̀2e���0g�l��ң�۠��v�͞3ώ<�[0�m>u�5��%�vBY�Qb�ΤI��fߍ�L�s>�G~jO����T�W�F��'�^olOM�\��R��c�WβN����r{�������k�c�=֞~�)��}���[�m7n�M�2������ic�������=k��H�Ɓ}��������ε��(Q�g�z�g�֬]$��n�^{��s���]����N=�e���������$9��6�7����:*�!��Y@�0��̙��l�p���^�,c������翴�~���2t���uЁ����2��>�=�H��J8�c��?\s[p�Luw��\78x����K�J����h�����oϜi~�B:l�h��������W} ��ζ���9�[dD��n�Սn� ?}�R妨�#���`���Y�pzu,�F��:�����̴���K�Eԥ��9i��Ni��T������ꭋ��
�c:�S6�B^2>c�/�z�)��n�����&���O�$��իsձ��'�\�|钣/^��O�Wc���5Lu����,OIM��p���:�R�.U�)A�2~��h�b¢���B\����Řy<��)����ϼ|u���ϗ"�{�[�4=�w���S���V��\���or/Wy��].�����s��}���{&t<�FII�?#ݢ�"O���%m�&�l]���gg)
D2���ufzVf���IMO���?=O�������*� MXfSsS^]}]ammM�ʕ+�%`���X�Q-p�v�a����C�E��!���HJL�"8�Q��	��0����R���·FN@H�.@� ��;:n��v���>�n� \�gt�Sֿ����|���%��u%�����.��b��D[�x�=��.��?�;����e{쾫�ӎ���O��j��=Ҫjj��s<�q����\nG~��3�])ƍm�&N�-n'm1�^y�u����}�]�\y�����Vەa�I9V+{�3%_8��?$EJfRZ��:5���>t6?F������ֺdpGV�@I�B(���C���.��Kﻕ��Y$)�2D��şC\������)������]I�F��.�	n\����e=ͪצ��,��;%_
���e�m��eV� #�;Se�b�wm]��,�L��i�tZ)�5�Kq�Py[TVѡ�����e8��˲ֺ�`�b �)$�F�t�It�<�&�kk�w��i�J���z(���[e�a�R�d��������ݳ�M��Sg/<��:IF�1_��Y��0
P�o|�A[�J��z�.#E>���tn�Y�UT����O?�w�y�,�/��u�E<����
g���3��(�s�α_��Wv�Ϳ��Q��|�bʖv����с���s��6����m_�g�UY,(s�Yr�2��Y�q�c���S�W��q����乆��]�����#�mñ��?Wy1P�R����#zg"zl��J�k����N����\�0�X�USS'��+
Ш����ěq&(lN��@��nW{)0��j0���g�F��j���u�Mu������L��	�r�e�5"����Z+�/%�CnSܐ�(/���d��
�75�h![���#x�T�Q�	�t��~݅��
3Yat��'�:"_�-�u������2?�ȣ��g��e>�5h�`�0~��!Y�f����"?m�tw�3flX"���L�c�=r�N��h�BcC���g?��?��+����I��rI@�U�^��82K�6�C��o|�X�m�UT����7e0p�5�����f�m��1�=q)���c������ϭ �PF�Z[�Z<�:^��¶�:���kO��_�p����;ݽ�>=��Ӎ�F wҧd���k�^{���d�L�����fN��v�!DxpTTT�r�,�Gi��m���?ĺa��g�yV�Z���YB�*���_y�Q[�`�,�|Ȭwyy���a���'����,k������Y�����C�r��qO��.�/���]|�g�Ș7n��G.?�~zٲ�.7p�C&I_�t�{�!�1�����ĉ,Gr�Aեm*�C|�d�u'�v5�j�J���cK�{��f���?�����;^����H\�i����ȡ��gx�>�1��,-
.�|�΄�F�vU�F'��w����D[�j��WxЄw��KX�E(W��g�0;'lm?i��m�-����։�����o��6��~�m�^�M𵇯H�u���{�׮]���~�%ttF0)�M�	�h4t��9G&��E���g$ԡ�	hNd�;���:C�Gُωcr�3�y��#�4I��(@p��[�G%� �� �
�yG:<#ߘ&�y��7�tyq��!�͓gt�O�V:���L�O�1jǷ4b�M�t��<?��5W�Gm�[��_K)A�B�3I����,';WC���=�����x���CǓ���z[�f��~���[o�E2��~�M�K��� �n��f��Ͽ��H��=��]݁��+�������γ�.����V�^��.**vZ��@)u��.;�3��C�_�ꗾ(��O>�p��#~�Y����e�FH�8��H���O��qP=�����-��h�6�ڒ�"Y��:j�l哓�l�>�r�r��t(>r�<��eG���{ҝ���37��AZ�r��4�hMΰ�d�ŗ�'e�+Iy��PBQ^���-E�x��0�$>�����ewX��a�#q������$vP���̬�"˾���<)=Y��&��C��i���lNf���P���-]
��?e��O�� HV;���d8+�R��nۋ�>�q���%�Pi���}kX>��ĐJK��ޫ�(�(ꢪ�D����#�Z����rӻlBy�U��-��MW��:�q�\���?�@�ӟ�d�Rv�Ͼ�-#�Mfw%� ���bیm�x�P���
�7�C��I��2�RFi(�s���}��Y��c�b���!Æ��_|n���o��f� �n)O��0ʉR�!��LK����(���W(J���)�G�R:6�'�=
�pEFJ �`�: �?�������+�F��$▕�wٓ,�5k��E>㔞�ً��x733M1�e�a�7`�Qv�g��~�qy��{���d֭A��F�ncǎ���J�����I��g�ң��b�K��<�Џ�.�����V��죏>t�>K
t̛+�L�s�!x�:E1��ҋ;
-q�*;���B�MZ,���={�������o���p�-6C�#x�PFOvn�� |�9Y�fn�|�w� Uꋙ0����/��O�/Р����a m���v�=�ڃ?��Thl>�l�P.�� �E�˦��U��zo'�DF_��0k�<;������3��J��v�A�|m�e[��x��
x)��6帠���juj��og���*�Y����l;숃$�jT��ɭgeHM񴚚Z�����3Oة��b��]{�ݙR��쨣��zP�8*_h�;�����?r�1�)W�^n��/��/���p���S�2��]�V�]d��v͵���ξP�RdH��I'�b/��ϰYB�d��v��e|;o��o����������`�^z��wٟ����� �F�p�M�����g���ku䱞3d��������7�|�����A�-dZ���/FF�ɞ��s>kG{��v�}O��}������Od�~b�V��*��I�����˕!U��v�ŗ۝w��3H�T��@��㤳�{�x����ǟx��V��Id5.�:,���pG�-�����%ea��X� k��c���i>��w��΅�f�C6c =pf�7�{���]y�]҃^��W�����s� � �o$���+�$r'N�أ|����5Uy�%,̲�Pn�YI˖-K���.;��V�^���¯;/7����3���*Y��Sʧ���̌����.��K��H��`⽎�����]�wKθ���*�'�gȌ$�+��H��{{Y���a��N��8X�|�����W5�Շo6b8�}� x8ح�]�ਜd)<�'������XoAg �8ć~�E��S��C�{�V���Ӌ�ipϕ{ �����8�8?��!�'���K�3����G|�4�#�AZ���& �!�4��5�x�9��6�lT0Z�O��E#=F_P8�QGߨp���.�Fmm�O�2:�.1˖,�b� ��shI��e����X��G�`'���9ۮ�pg7 ��w��W X�n���RÌ�:]���o��V���� ��_�l�6�����{�������ٝ��t�T�x�/��K.u��K/���K1}��'��뮷Y_|b�R^3�qO��������cOX�:�K/��!����,{�d�2�R�
-���R�ڛ�,K�j��ٌ�/�qa)���2$b�&l\��$^���1�!��꛼��P!�AJpS���\K��"����]10c1~0p�c�������8otK!A��b�!��2����j)% C�)�XO�^��Ьd��&n�ɖ�%c/�Gf��Bs�5*����O[k�uʸ_2ہr���n���Z���6�jkU���e��Y�*��g�!z�v)Y�87"�dl�(.�^OR��ޙa��m7�G8$��)Y4�����j2>p?,�N�~=km�7Y��Y>�@���V�@:����d�J��ŗ_�c�>�e�w�3@^�m�{�/�S���5p+�A@�� B�piT��}� 3Kh!�&E��h�~�%FT������Y�� e�zV�e�]�̠���>Q���.�	w�f���er��3fp�m�e����pz�<`Ƙ3g��~;W��|�u�GTqc�Y3���"�XZZ��e�]�M#�{�CѦEe�wZ2��Hwnn���A���������A�0�5�	��z9��`�)����Qb\�&NkS����/\�k\����bu��>����� �>������e�hǝf8Ο|��čy�K���L�6��6Z4_�V�@b���H.s���J�t`��w)FRஶwd ���	F���F�cխ�*f�p+��B;�`�`(��޻������*#Q�ݐU<hG?A[ 7���������b�.�5kW����B9��~$�AB_�^)H������~�n ���s�{�d}�T���b�!M)7�&���xxC w�jݚ*�x�=�ԣn -[��N=��v˯c�i��&��,���_tl��CI��g��m��V.�8�����}�i�(��RAA�r�a��C7��W��u�*e�}�.����UU��$.��9��]�v6}x������b���f�\s��}�z�bJ��O��ޜ�/�km��!v�ǺkMM�����8��F�AeX�r�+�l���t����:����v�u/�ƌ�o{�]q��aU6rt�]w�v�aG{"����8k��v�O������-�q��L�(�r�+��y�噾�+�.Ynˤ7��l���m@��2W؇����1G�-Q���c�;�~{��d��}�}������3��<d��S�3�<�n�Q����h�@���+|�\��e$<�w�Z�1i�cȏ(�hWĥ�Fm�oi'd�8^�c&�5��i��-�9_n��9�mÆ������/�
����O���X�v�~�[г�u����	�dp�=���5�*S�dU��|�����ޞ&�+Ye�hjV�4455gI�@��=�uY�aԮ|�WͶ1_t� ���<K�[��z�ʕ��E�_w��w�N��>)�ݭ4�D��eee�D�����VZj���N��K�1�:u�PY;��
�%G[��M�mʔ�af���-`��Ӆc��K�l�����?�����K���;0�1|��C��f4�Q	��:j*L��gB�o�Y�C��Q̹�@�����{��q� H���A02�<���0,�����y�o�{~�qH�+���]�	�qF�H���'�Sv� ��A^�㞼xGGΔ4�t|>"'%�w>�#��%_h�sv1���!��/�r���&�Z�4L�=|�ٱ��$��;
�1�÷�	�|��IR��/Æ��.��]�~z��/�7�����Ův��aS���5 �	e����vʩ��C<`W]}��擪�[T����w�u�a���n�ɕ	���n�������撋.���F��G�`�
�ϗ�m��Y�:�C�Ǿs��&s����j�Pa%��Yr�pK�a��KP��Y�h��z�L)����$�R3�U�(�2o:��~�T�԰�,U
��7 ���,)��^9��,	kh�.%��"�!E�Rw�3���@q���)m��I�f���V��O��
2��"�p�9������nkSٓ�n&|����r,c�0�dj[m���e]AO��gg���0a}����KV9ը�MFPc�ґa���g���I���:(�ʒ��am�c~C�N�[��์}�q�+��N��L�{����8Rz-2�S;��㶳W��K�ݏ����b�mt�:�:�K���N<��ns��("��kx��c�C6�>�2$�$������3�cL�.e�tP��rC�E\.�/�I�DfF�'���0��L!���;��0��9r���Ϟ$Wpki�$��=ϐ�����QF�5�o�<6�<"�ʄ����r��k�8�a79��q����]H)Y�~��ն�(�,{�W���.l� 
�����)�+�1�����Z��E�9C����w��BWWd�ϕz>�!��@�8ֶ���͙;�>�R
 B�1�Kf6���]#�-�Y�A٩ӕ+W��k�:CQ�n�c��W h\&�b`�@��d픰���.J|d'u�J]�+f�R%_��V�7����_���9چ�=(��E?�+�?��;y���8����,k/�s�r@X�շQ��C��l�h��u��O�|����w�{�)eE��@r׼��w1�Î;�`{��3HG��ڠ�}��	��a�}�������5���_ �Ȋ�k�nH}�A�͵�b�*;�����~�23�l�|����OKo�fl�>a�͓���ܨ6F�K�����s|���ǎ��kVڠrf�F�U��ʿU�oJ��_�ǟ|T<�Ζ,]j^��^)� =���v�E[E�R��V�����]��^��N������w�F'��u�m�i[�q���[#���~�����G� *F!2���y�YFXQq��s�m���;�H
��A����l]�*�0i�]��l����d*+��SN�g�}F��a2�Ǻ���;F:	2:���x;b���f[�:�H�X[e�U��NW��;;z�߭kY!#{�}����f�*���}�?�a�����x=����"O��P�CV��s�y��9��eev����p1C�����H{�m�I팴�����Fh/�Z��e�x��h��9����~�wY"y7f���e�2��,�$gˉ��������l��Ş�?���zfȭ���=}����֖�����$v��G���=�]2J1�Rrr�Sdxt�����I]��l#]������n�'�G"55M��� �|�Q�V�t)}�$��}NVv{gG{w}}��kH-� �c�6��.˙E��֟�~�޵�w��u��ݢu���$��U&YgJj�T������
��j��E�%�q�i�*v�}� �������|1k��ꪪ�҇G��וʊ˔��P�U*��{��Z�l�ԩ��a`@�P��
ժP!�5�������q�0.�0L�E&&>����=W��0#��4T���[��/2,#PX��^0-��JzX�(t�.�2��L�b`��s�GF��r� �}Fbt��hߐ6���N��i �����7��f�`:nN��=_e�e�Uⴵ��ӽu����*P�H��夌���`W�P�p�&����E�>3�Ko�AOҢ>��k�O��=��w��%�q�?�A��>I���#����v���H ~�^~�;�<�w8�#��w�}�� ���G uςH�a-U\��x����[�?�k�_q�m������������vr����uL�SH��T���qC���;���wb����I��m��~6n���G�p�Y+cl���:){���:kli���&7�*E�uԟ:����:�URz�QhS&���S
l���aJ�m;��fl^d�N)����o�lQb�
��$�~;j��7���d�bd��y��y��Wh�ϲ�fȘKW�=V��hmMV�Tm-��,7��F���tś1.�v��i;Mɵ�rl̐,�P�5�Zi]UՖ��`�5��Rg�ʳm�-�l��6j��lnEj���#c�E��;ٚթ�\We��Kk��u�7h�F�Fuޠr�H�d&�AiWV���ѫ��Z���|)���f�J[�����Ze6v4[[O�ȲAC�E�����D���;��ѕw�2A�����d�y<� �aC�3�6�*�"k�5mq�x�S)�(�,�� �0Exx	��E��y.�/�W���k�+�X�8R��ҿ6��, ���txNڴq�I� !����	���c����BX�R�q���A�!M��B�t����%/f/�!%/OG4�Ø���x}ec�*��\���0̸ϕ���L1[�������O���]aE6�C��Oq��RD�"�G�鮔̾�y!����c�LF7}|Q�v����x]����蝤M��!�����(����=����5����2����F}�|I%�~�%f�5��~�w�1ec0�r�G��	��P� |).r\eq���{� Йs����] ϡ��;��$~�|b ȋ��?I���!�>�$���Cf�๦f�U�O���aC���f��pc�Q���sP(��ۈ3r���z��x�x{����pX#L]�&�5f�����k��hx��(�d���ם������D`P�]�1�?E�G����1��|_�z�Ϩx�6E�9<RT�g�Ok�컋������sO�A{��ر����0���a 1'/�;f0΢-�8���.����7E;�և��û���^8����Q�|�	1�F[��p�..��w<x�;��^�[�z'��>B|�ġ-Ӷ��Q�i��8��{�`�UVUe��e%�w�'�-�|�yٹ���Μ���.5]}Q�ʘ.V�Mb��#+M�O���O�<d�e�����_�,��ZPP��H�99�,��7"����6W�Z�$�Y����,����ɠ����}Sڿ�ɖ����,5rt������0(oȐ!�
y�旖���,.*���;L���ä���;|ժ�#��]�f�D�fꪕ���;w�ޟ��Q�g�>S2�O?����z�W�=�ܾ�Օ%������s+�۳��S����w�}���������	}��1o���	/���w����~����r�w\����n�?|?,�� �b ���E���>�+Z�Dt�b�u����Y�:���TH�QhPhTA׮]�(��QFB��kt_�d����3�,�=�W�:1k]źuuʯV�ת!��Z�|j���{�Z-��#�6��G84��tmP|�5����Rz�S�6(~��BL�N�['��R�V»YL֦�ۅW��#�ub����r]�)�R�L��
��JaA��U�u�nmo��X�B�{��YR]S�l���˅�2}�X�����U�����05%mqWg�R)X�e寕�TSQQ��av�QIa����!`��	!(h�A>���4V�2�A�"�$4z:K:�NT��M�4v����o:���c��]Tnϓ��C�D�D�cR�=o�"�%|}�17�X���@��z��PH# ����_�]�c{s�;^�Çڀ�%�&r�Yg�5��Ķ�nG�6]V]S�(�2��)C8E���ʵa���Pu��z�d�{�շ쉿�͞z�E����_Q��30}#����"qh�tƾ�����T:>�K�R���ck�Tج�����+�O���Vk�Zg�5Ֆ��l���&銥¢�
Kҥ��Jm����_,������k�,��-�{�Y��c�o�}�pk�ჳm��"?4�JҺ�<7�v��s���4S��Ym%��,�(O����s�l���������~�#ڿ��{���O�~m�z�v�Rg3HT�2K��8'�uDt�����v�O;T���m���0r%dJY>�L��Xqn�u�����e]28�,5S�URl���S{��W���^���4#ЁↇK������oӑ����y:�z�����l��WV�]u���Tw�c16���A�ƅ�E�i�͎� �ұ�BGJ�1_p�v̐�����Z��R �Q��mlg�l_�� (�4��PVu�{�$u�>sƳ�t��+��+���������e����b�!SBY�)�OG }�|��8В �;�!�S��]�2$�
��(��cź
cp\�0�Hӕ5}"��x�-�c�ex��1WX{i�7<c�!W(5l������s���W�WP�p!��#P�W��G~ �&-��"�:d��A��q��ɕE��vd%x��W_D��#m���A��S�	rz����s�� #C�-�W���e�u���cp!@31Q�	�C"DZ�3 O�HA;�<�R�6�3B��0C��ŋ��-���=Gq�}��oy�.��7�on��|��[`�>rÀA��$٠lЗ�?�Ϩu�s�)�<��8��V�#wC�'�W^�o�|�[0��=�Y̶�Nw� N�퇴���=�w�f���y@vL-\h;ﲭ��VVR�g�8�z��f�֓����/�����;����o�͙{�����Z�F�A~���Pf�1�H��S�.�N��B`S�♂N#��񈴠��6�' ��7y1P�w���܏�cd�f_�o�=���)twK���m��E��� ��B�b�"���<�la�WD�x!縆u\\I#ּ�g�=���$��!�3��������υ� Tp���P��,�EV$��_p������bכ��tb��n����p���U7�ˏT�m���o���Az��F�X�|i����מ���!]rpfzf��/�,)�藕�=T�v���~����
a|�h�?�pIeE��ʊ���J��:�,	��j���T>h�:�䶎�<	�\1* �)H	�Y�5b�ukו�S��V�R?ҝ�h�%v�ʶޝɩ)��L��[{�/�R��7]�����CB$]xa���2^�;��0���3M�+S��&BԪ�+n��&�t)�%J'_�g��m��Y�P���qT@�rR��H������S�{���W��fJG[���T��$$�$w���u� ��H�KR��.ᔫo
��0����J'�th���0�=�D�P�(=������%,(���O�sN�?m���^���;0�C@h (.v�C���&����]l���^���~��[�:�{��G;��S=�p��l]e�FD������|w�7^{��W^i�]v�/�]�j��u�Y��c��*#���f{춫�������;O�D��*e{��n��}W��2����_�M�0�z�o���ϲq�ُ~�C��"{����Y5�;x�5��e 44��ٳ>� ����Uֹ��l]�e��m�߆�c�$L��p��c�8A��nф. Y�����R Q��Ӓ,���j�[l��/Z��9�o`�;��ՉrХ��bɵV�Xm��96u߽l�6|�P[e��y�{�o�[kC����r>l��!���U�*X\�m�G�YGs�-�|�-x�c�YeӦ�1Ub/��U�g����|�/\���[Y�"�P�ը�^~�9[��'2p�`+-+�\	�!���	��R>;dp�Z����渄T��)z�UwI]RrE��B���QVTj��ėumR��ڥ�*�+j�/�'O�e�Ջ��������l���|@n᜷`�z�a�>��Fb;!��zۭը�C�dM��{�i���g�Ӈ׮]����"t�O?���'iR[c�r;F@l��]-j}m�@~@lWN2���?#1��2}k��mn���|K;�1��O>ț��t����弬l��b��a:�쬰�eȐA~�f�jW�p���4i�m>u)K���)mT2p���T��FH�C�e�8�|�+�d��&��鰉�yOqw���ç�eko}�؄��U8V�\)R�8ׇ��t'�+(��Ց�%��� 0n��a<P>F�i��N�p�����h��QGaL
���0�^��k���BT��p��v�O�_��+������g��kXKx;��;;���#�(�:�k��GG�O�:���r�2-̢�` �raHQ߮]4��O\�!oq�{]/_���������7��Cl���u�2����x˾q�1VYUa�y6i�;���\A�v��z��Da7���h�nM�����{ﴏ?���{V�kj*3_�6��Uv�A�ښ���M��I��{�}���NNJ��}�l����ڮ��l'�x�}��o�ghc���:{�g��[o�?z�w����q����k�����K.���f��Zw	��9��Sm����o}�f��������b���q{;��sl뭶��}n��@CPq��x�](�ΙoS��d7��z���6!BO��y�}v���^��c|�Νw�ӓX����S����ϫ��u���������Ɓ���D`���+V�w���1�e�<"{�q�q2Zsm�*�����ſ�ǣ\��`�a�������������]�LA��� �1�v�E���iS ϸ�� �m���;�Q�1�(�b�ev�����v���SO;��믻����)m~�᪇�%��QY8[�������Q�F\�l���q#�\c�t%>|)�]�	���_� ��ȋ���M�/4��\��p��QO踒cU'�p����ϯ��r�I���V���^XK�)�����o#^���A�g̜�v:(|
Q��s#-7/������>�����/8"	��r��U+W�VV�+\�di�:��A��������ep��a����b�.��U��#�:�2�	�H�Ҩ�Y�d0<:e-���K�� �}�$�S���"�S�t��s��,�I�%�o�/�l�@~��ݔ.f��ɪ��n��>b �{6�U�O���w�a�}�YobZ�WB�p�Y�݊ӟ�c䡡����8�����etF�A6����?g�"�,�t)t(8t�o7C߬�E�(Dt\���4I���J���~���+�P��S�f}a�_~���e������Ÿ��w����曻���v��LO�_~��/�\��|�A�@4�̺����o�ɖ,^d�&O��F�l���>�_��7vх�f�������5�׊�����-���N;�t�s��lѲ
;�ȣ���F��&�Jͳ���^^�ay��Z�f[�F
�}dUkWZq^˷BkZ]e�+�X�ʚ:����f++,�gm�d�8H�Rev����JG�@����f	�R�V-��%�kV�N�DO	��~�%��������5RhZ���j�|�0�����Y�x��^��ꖯ�N�]鷫�>e��(���56�_�m;}�:�v��Ŷ|�Z�]�d��YҺ�2b,9��Zj�-)��re�1�&n��er�x`�:���z[��lU͖��� b})|��+��Q})���w�KIN�)�l��!tUf�BWo��2 ��):��Κk���7��ƨ,���>{�-�/3#ݦ�ok>x���Wk_���7UX����V)�������=�̙��;�p?(v��(й·�[/o���N�xp�]yՕ2��o~�[�`/��b�I飽p.	��ߟ�G��Zd����,y1�G�ͭu蝮��Y+��p�}�q�<��e�W?��TK[���x���ٲ��e��X^fQ@t�Ō+���R�j�
/omM����C��mP�qo�̠3f�����?�E��a�-2dt��Q7Օ���xQt~c�QvDc��x�����5�8F-9�l��Ѣe��(�͆j78۬K�r�uD��C���� 4@˿����q#���T��K#�(W�)���7 e@)b� i|ed/H����s����d3�ʉB���>����y��7��ok;�>��(��"�<C�:ux�O�`,�~���߱�
۰����_#�����!o����RN�0���W��C��&��\���n[7�)��w��uVE����6	��8) ��N4�(��;���"p�G�׬
;�-X8ǖ,](����O9�w�KO�I�Y��T����Z3Wu�c�GO����8��������?�*�c�p�3��C�k��=>x��@�A����ۢ�_RR}Y���UՕ�d�[�h���Y��_'Za|%�#���;�|ѯђRZ��8�܋�.Ŗ.Y�~�۾�!�1lH���Iv�!������A�f�F�	`�A3�F�O�~����?�f�W�U�:�n����63�V�������ӏ��z�ݶ����m9*H_|�����«Vm��~�ӟ���Ȧ�99�I�LF�UW]e<�g�@�w�qvӍ��~%���
;��s�G���	�{�������j���%�/����������9������Z�|R8�C8��Qf��H^#x]П�<����{���۾�����d <C�Ef�3����g��~�m�]7x��>����������#����������i� �}�+y#��q�Au�.���q�W�c���E\c�>���b�HPv��Y������zF�@3pm:*�#��q��C$��%�8��:X�d	߷L�:u��ѣ����U�UJk�p �������]}�t�}��Y�K9������ȟz�:L��̙3�I6]v�]��ՑN��ִ	���*+��?{���_'�lWul����0���l0��ҹR��8
S�8��7�����2�;P� \����C�Hr!0j��1lx�I筷ޔP_lW_s������S�<c�}�7 �b>䠃֋D�4�����v��������������#w�~�d�٧��+���K��o�c�9F��?��������o���Km���v�}�˾�m7u�]q�lyM�=�ڧ�ym���l=Ń���s����J
Kmp�pد�:�д5U�ʚ*[!�[&�@KV�� ����n�'��f��#Q��ҋ��3d��g꿱i���%[Q~�-������Z��U2�D�6)\=���m=Ŷ�y+[�b�-�������E�HV���f2���G����ڬ;��*V/�iSF�1G���>\eO=:ǲ���;I�E�1}�ᖙ�`s>�k�?Zd�5�]]c%[oa�_|�ը���l)�G)$R�Gn6��e���G�����VW�Lm�o�mm�^{X���:)���F�P�N`�_��~H�\��d�iqn�-�o���-�"7h�f�ٔ	�&�S�%��NMI��cFZ��w����9��ł�` U�[a�H��@�� �y��E2h����4i 0m>'��8Q0��\sό. (Ќ�#Xq�@q?n�:�:{���d�/��!EN�D�gg86�(�_�)¿� ��?�;�:'�>�����WM:�cԏ�f����"�Ʉ�v!D�2�ߤ��;0�:Q��Ḁl_��,Rt�cf�X����O>!HƉ�_�o��N��:Bcp� /pEi�<~	n��� p�S�CW tiB�q����t���w����b9�Uc�M�8�?�y�tЗz��П���{����|�aJR��1����Ί�/� i|dZ?�(�l*��N��)�|_YU�	����:��3<.��9��٥k��w�[o��h���.x��&��9F �j�	=p�����,�����v���+�o���h�l[L�B�&ٛ�gm֮��(�Z*e��xx�$�>x����c�g�b���$�+GD��~��Zh�r̛7�f츃=�l�x���yR�Op�{��fX^n�UT��ys�9���>� ���yz--�\�{\ iԥG���<=k��h����8�#}�s�Y�-�Qq�-X��l�}���������@f�=�{v�oe[n9��K�O�o.���>8�Z4O�0�@}G�o�jה��p��%K����lCΠ��I�ͳ����o?��U*s0����c��c�/�����|��Kr�M#M�TRwR���*P�P�²��wX�x��HiK=uM%������.��s�=ɧ�������ܜ�ߟ����̙�3sd�Go�U���X�����	��M^�m���v���{�=��OS���j�AG=���p�1�\|0Frz�|.چs՘Q�;�N����'|Y8�ܭ#+��ۿg'�p�ʕd]�v�m_�o��*f��;r�}�_�#�Ā2۽k��x����W}�96��_߶�����3P�C� Cy�W(�A ���~�����n�e�7��F��׾fyR��U�[n�����:/!C�Ϩ�P?t��}�?>-c�#����~����a�%��'��������f0 ��>,�ʀC�: K���{�M��`݅� �%+�"��O��W��>j�w�������g!��w������%��E�VPy������/�ï��D�{O�Hz�(p�7X�������:G /O[ �<�2�?�D#���� ��K:�H!�����C��@R�����<���菩?�!K�rfmUS]�V�.�� ���=+� ����<Ҷ��������)�Ħ��i�^uջo��x��5�x�)��n���>�!��Gyd���s��P�]��`�a����<,�C9@X�\Adt�t��?�E�o�.E�)'n'v�d�g��u6�r2:�{Ա����}���c�qE��)-�&}�_w�E�M��\�>�)R����R��4Yf��JGʨ7�s��T?�p;�Ӎ����\$�a�y���'������y�J�w��v�QGپ�[�y��[��f�2O�IA�����[8L�J���\+Vj�CK�C�����ԇ��8�Q������
N�pƑȔNuhev�񣭬0϶m��=�wX����:��*T��[���+�X�>)9Y���ec&�ک'���ԑ�ۦ-����d�R�zd|�'�rճ���ƍ��k��4�f�/���R�[��9�[x�3�*��Z��vm�e�C��X���3�9��,ȷΤl�i�Iδ~F�ˊ-K�ro�%)f���<$a�;i8n����cG��>h&#9��J�����a�S��N��	�������\�۶�\b�ʋnѱZF/Q8p3�f�:)@wy:t�@�؂�4�=������(����I�(�,AB�b$��(K� �5���u���2��������g,C;唓�4�%�GPx)|��w�*?�����EE�n͑��1��7 ���H̐@����P��x�=�<�?v~N��"��������	tD,Qcoˤ���H
$���`����{,�!�M[�J��󴙵��t�a�!Fy�y��w�<� :F��6q����{6i��{��d�0K��M�6fФ�(�q��7dm���H3���]�	3�7>�C}1I����A�A.�4E����*t��\�`8����:c7̄c7@	�E�3�&F,J?��8"`��e�ʫ�8��&����ݹs�V��hvÀ�Q�1Zq|�Ql֬Y6���v��y6q�x;n᱾�x��Y6s�?c��s϶#�͔,�0tΕ�ex�"L�6զN�"��(/�c�=�y����?��	o�%�����=��]z�e������I�K�xk��Ā[�d�h�0��_>�5��3��ĳ�C�w��<i��c_�*��tfϞ�:����3x�]wY]CXJ��Cf��}7�
�{���|��6Q}{���;�c ��9�s��gZ�J۳w�mܴ����e3�@��� /�}*4R�w��rډ�s�l����x��3��7������� wu��3�>g�wl׻<�f�Bʠ��W�ԯ=��3V)|-yi�=���6���_p���חڋ/�dK_�3xv�p�3�/˄�WW9-^t����I������(��K��l���]cSnf�~�������t�+�a�K�ʴ�j�{����[��浶u�&��N����up��g�w�Ɠ��x���@�=��Siwz�g�)`x465��/�իV;]Bw�(�:���*$�2}�w"��k�6��B�D���]>��@y���%�ߓJ;��FY����'�G����Q\o����<]�l9�s���n����>���'�<[2q���d���J�U��`��~�z���X6� <������k �X� ���z�]̃{�-��ߑ�`roLW��<����Y��~P�������aKCCC�������鶙�o:��l]vf΁r�^�/�����B��-��O�X�b�� oH�d�|%Ik�믿~�:��Q�GY�$4Qrxt�#(�z?8�� �`��g�|S\�>�DF����LU�%�7���M��N�0��(J�v@�����<`d�er)J%���n���/,K�DX#�8s��e�j�j�F�A�gԎF��}�<��>��#>�J�� ���R)=�Ԏ��O<i_����W^Qy{m��Y3gۮ�[�y��gUXjn�u��Q2�U/�գ�W�UZ}s�ed���d��\���r,	<���21��
]�B�gS&�l}��s[m�k�y�~��o�%�V0f��:�F��d���[eؾݒ:�l�IJKon�-�Yne��꠻l��<<�)������Pg���ky�6��b��������sӥL�#+��q��P�Q�:��|�)\��m�ܢa����w�:N^o�Ϸ�!�m��V(�&e[?k�{:,��,���U��1l���%�=EW�I~b�����}S�%V(��}2L�gT�����Zk�r�
Kj����v7���jjl�a#�����U��8����)
> ���#Mc 1���ݢt�ԠĲQß�Y�7�r<��C��z�Z�l9��V���9�c��3O�)�(U�2��1��C�><������_b�����߮���~F�1�c\x����R���F�g:v��l-x�X����zr�w�h���{�qe�3��a�@����eC>Gi�U�Dx6*+ �م�?t�1P�R�(k�K��s��v"=���#΍�a��P�+��ʞ�J3K�srd�3��i�9�j'�ic�A;�	���5�`Q�ٰM�'�*�#�<� "���B���N��o�K�SJ=a^�Kydp�b����w��`�|��Sޔ�S,Kt^UU��b��.�p�y��g��^�0����I��{~3���;rh��ufq���6���e�b�m2>8�8S�l��d���v�� \��!@�B�s��p��嗽� O�H��?ھʝ���z�>�y��O�b r��('�Š|���}���k�����B��W�C��'�1� s�m��4گ~�k������=R��b�D�`���o�;[�v�ϼPң�0�0h�Kf��0��=�SkDU�_m]��􂢏GZ���M���ē����;l��*[&�,/?�JJ�mF�̹Bq���.[���d�gMK�E��VRVj��L���ْ,k�dᅁO�eS>�+{[�F���*۹k�x�_}�0�(��/��76@����^~�%���p���SO�]��w�x��^p��ؒ���'�x�b�=�����*[�r�������_���T����^tϴ̰=�����3ϊ�Rx���OƹV��|�93Hx}����b}C���d`mt����>�G���g�6�x#7���}����.�G|ژ��{���.��˫�@���(%�ʲ�u|���AD�]�i���>����󟿥��O:��'��X�g��6u|C��ee��@�����y��	/������8L������4�==�YA��t�#~#/i?�N����ч)
�Y��,���J7�S���P�!C־��+K���/�h�m�>��O<��c�.]z���d��0�H�@��!?M  H32@(@$\����� q�'B|� z���+g�M�r"F�$�~�G�*��� 6Hɣ�í7��?�яԙt�q�C�p�uk׹pcԋ%�?����O��?����>����=Y��j�j[�f�=/!����ؽ�?h?��Om��˰A,=;�f6�Ǝg�����]ՖV<��R��79��dX%��Xo7�7{���J�u�Ӧ��a%֮N�Sʻ0�#��#)%B��0�.�	!�𶘗�7X;~�p7^xv�-}e��ִ��X��	6i��4g��W C&˺�q�񿵹Q�E��6R���i�-3�g�m˦f۳��zաwlL�y�l�0c��H���\)-��-�ᵕ�e�:kh���l�J�	�d�gT���LO�:洜L�;�敥��ˬ�5��F�Q�����c�(��C[����|}�hč��K��8|�� =��F�e4�Cnq� �Yeϗ!ľ���N�o
�rT�nk��f��U���f�,㒲��`��O�%J٢���`�Nڇ7��F^!��e��#�m�f�v���f�d�N�r��(�#�%��)�R�G��6m����d�٘�����+��.ea�+Ot�c䉲M9.~��v��/Z��v�Ǐ�ѣFڴ��l����M�Ï<j{v��P�˹Pz@�/_�Q�YF[��S���������|	n�K�8눎���qC�#b,P^ E�������LmF�\G|'�% �Ep�e�e&߱g��5�=�� B�'�$�[���D����p	��=&ym���x���{��I��(O^�&�NG�S�A�-�K����Q�D���yS�)��H��q��qa�̲�/��N?�to��,�K/�T�s�/��8��k��h7�(+��2��QN׮[e�8��alt�R���G������K�6n��3
(�x�kQ[�[��?��V�\�W�M�ȇ�A�=�S"�,$I2�E�c��K/���,����yw�xڄ^=�=EKs���<i��z�f_��>�%(�<�2qoed5�#�#@UU��_���wL�c]x�E>��T׫��GF�v���oQ���Ax O������3�J{et�ɲF��-�Z�F����('3��ܱ�v6oܮ~�Y)�5��K�f�<��A���?�g�V�f=��F�;w��;�[����lھ�V�^�~v��a�I`�����R6f���������6w}.���_�gg�y���x�?I���Ջ��.�c��|��G���M��۸i�����W�~[|��:D29����c0R>����c��)�J38��tf7����9�g�� �p0v֭[�m����7�<�'=��I��e��w�6��op't��m�=����(�1����{_6x���[�V�� �K����ؾ3�<s����O�f͚=��瞿����T
8�p���!W~'�����P
�&�?��w���~3x�����@��T������`ɢo �TQ���� �;�#?�Sr����h��g������Ad޼�o��3� I�Ї>����ǟ5jT
�\g�:26��!�H NT0���og|W�!� %6l��9ip��2��x��ѳ_��vH��D�%a�����n��&_�����%�y�ط�w�eFUQ��w�Jz�(�XB����A����7�T&gxnC:(�|O��!a��P'"�ѥ��B�@��n�����ԓO����k,e�B�ϯ���b)�ɶu�J%-�2�2S�H�-,�%['�ΐ�d�[J�E�7��l�^�㸴��{��>+�˵�eE�~�[�z����V<���5�ʇ�PL�QE��Y~8`Uum[�@kS��v��uzY���/#��3�R�2eԵ�.)H�9v�g��#�m�F۾n�e��{7�X����uV0k��s�Y�S�d�������zSm���c�>[�f��Zs�nkX�NZq�9�X;�����^������vk>S�S�1@7(���d�p0�>Е�Q�4A�%�5Jf{_�eK��_b+_z�vJI�t�1o�p�aՕ�*%O�=��Њzl߫�؎W����ꐋ��C�k�;�s|�݀_��.�����6PrP� �Z��X��2+D��T���#F��3g�⅒<�uZWt���n⻺:���f���6b�ߗ7f�8��އ\1�P�Dc�	Ŏ�Y�f��y���}���x�R�pp�~�믻Q��61J}/�<������L7��ءy ^#���*3��{��C�fO2���+�=�C)���ɒ�j4�\	R\���d� ���D9B;�x*	o�>ʯ���O�D9�J�eyYyy�;�ٷo��,���e�g�[F+��(�ž|��w�>��ʗ%J�]iwZ$opȬ1���
�g�{�XbH@>Q��L���\�NP����0CD��Z1Ì�$�v��,��ȑ#�K_���8�Z�=K,�R�ժ�7�)��,�bĝ�d�q���v�ݿT�����W�ݻ���M�?㰙��̒�\��c�ad�~(�ԅ|iS��������
�`[%�b`�x{vmwϒ�#e�"���i͚u�$K�`Dz��4Cz�'A��:(��Q���Z��0p��AG]N:�$�= V�\gg�{��J둲��A,?~"IIo��</C��,��ho�EHK�p��#(��4hRe����[�� m�L���N��jS��O~�K����z�Zԏf�G>r�}�C[�<�����O�@+I2�s�|�0Nj���}�2���L���;��l+�As�)��p��1x�8guĤ�����N9�tɏ,���������~��z2 �;�hnl�o|�;
�tc*�0���7S|�!����z��s���V�#��<��>̗V��dq˦M2*3�3���{��ƨ߃>d����>�bV� �>�˸�4��þ��g?���Z1k6j�h�Y��я�oT��a��#@/ݽ�{�Ű�|�O�F|0��z�,�'.�D���]���5.�ٳ��0?�ɟ���"cP���嗽����wO�6�$���!���K�$�3��^��M'B�?@~��/���9~���4]]��<�2���c4�{�x{�9<�C�^��m4�����ק|�jժ]�f������9rPY���m�?	ǔ�o������'_Tǝ�����a6��&y���$�"�)��y�3���	�E��x 7���8N�3���w�T���������˯�j_t������a¾�(�(@�@�������g��
k��cP�N�RPD�y�Dp�(���Ѥ�e��r����f�T)3�K/c�E�{�[��sa�KY�א��m��l�Zu�����g[��J%�D���?�ʈ��L���hiyq�5��-�g�{�J�*���N9s�M�Rn�����њw:�Mj���ڔ�6�(�{h��^Ϟ�t+,͵)��[�ڤ����@�-j']~�M�UfK��l[�쑒�n5�2{�m��l3��3�J�$��M��bS��w؈a�a�f[�v�{��n���2��T؈�3m��b�jb4�Ҫڛ�OJ�@�p���:g�Q����/���R�ߊ����RiN���-��|��JI��}�12��l���@��-M8��f�����?�i����Hs�V�o��w�>�)~����}�{��-� (��Q"�((T(Zr !�_{�U��i�����;�\WJ��DIad:���m������묹�چ/�������a#퇷���"O�7��A��f��ec�-���s���VU�s�����QhU6�b�/�	g��;?�w��e�S��u��(���3���&X�^Y:ˌK�0�xO< �4(7�-C!.e ]p\x�Z@�� �:$�D��tȇv�r��ޗ��@.s�Qnd�F���6a�8�;�H���˯XZ�Yh�����裋�^0�(G�>Efp�h��8lvgc<�,Kc9��*K~���bO%�:�$̙0����Q��4i��~6���
��g�u�ރ�0���Yrf�ٻ���|G
c�}�k_�����X������2`v�wܡ�JqŒ:0��:x�83V%%a6 ��Y3��U�gx7ԏ:�\��ڔ��`�2�@���,'�}{v�;���%@K��;{��>�P�P��Wԑ2�_�����b:�2e��[>���MI���Y��Q�)���g��u	�2�]:�랶�G�?����W��-���v��N������'>���;p]_W�H}0�1��R���n˖�a�#xf���΃k�Il�h'��͸�.FfNn��ZQa��eXow����/ؗ�|���z��/E���3J͞~������α�Ņ�<4;�=�8�����["_2��ً�ހ<h�=>�N4ҫ�|���Z��s�;�]�3�J�Ҧ�=���z��m�n@źP?�#�0y�{o��;�Ӗ/_�T
�U����~E�H��� /Ow��f��}�&/��\
��9 ǳ�Q'����
��H�����I����(��{Q|��SN9���� �Ci�_w�/���M�8���	M�LB"$����;��t���	���~x�]�M���?4Pn��~�|��v�@����ia`�ҥ��=��O�}�ݿ�	�^�) ?�~^L�@�qa	�~�9@ Q����F�7˥�"�Qrtv
�@L�O^���tA���=E:w/砕����Њ��=6���BΥ���6�#�}�������9�#�%�Q�2ץ4H���T��!O�����s=�8���]A�P[K�+�Rٌ���kOc�Um�i[���������{l��[��*5�ғg��<���`�vO_��<^��U\	ց���d��m���Κ�/C���
���yv�$+�k�'�'��w�dO��;{��W-+gi�wO��V�����[g��I6|H�e�Iql����:\oY�P���<۳�ٶ�Yk{7��w�{�8�׏c�=�^z`���ه�?���v�YIq�{`ڸz����e_�eu����d��̉6��[�������ʗ�� PG��m2����T���*�/t"µ#�+�_�Q��W�-2�L��
�����,㭥�v�Zg��.�>�!t�R�n�1���56ݓ����1�(� U:�Q���7��wT�GI�bp�ϙ�j2�i�F���ֻ^�o���8�����X���Yuhi���|���]�Y�+c�]js��vc�Y��<��7f3pMˠ3ԉ{��0�bA�^��C�zx��I�ub�\���f� o����%�����2 x!3��2d�7q	�|θ�e���Ef���DQ6%�!��A�g�)7�@1�ƈ�l:ߡȑ�ɐ�H�X��y�=��	K-��=�$.������ >&_~S�X/څ���&�`hM�Q{�T�8O��&63c���:)���D�I]0Z��á�0�G�c#�g�l"�a��6b��5s��)V��!�-.#9G
�����gۘ�dfd��n2P@����Lf�1�"$�#Wp�J���à�|�t�W��?3������`f,*���m[|v:�I�3�� �
�>�g�!H���=�YpWbxP_��|��@7���Yg:��F�Y�͠O�Lc��i'�a�'��2���c�l[ <��6w�L�6u���x�{��v≒�'��;Ǝ>f�-8z��?�;r��7_���Qz�o�s�yP'N�Ғ�*/�P��&�ښ�۬��H�b��/�*Z���[>d���W�_>�Q Cm����%�{�l����}74��d�:3x�y�f��%/��x����[o�o��F
�g(2 ����|p
��3���?�.��c�2�dK���wEٝ������H��	�p�e�V8 >���Q�0Ѕn�1�� ���\����4������Cf��e�}L�����LVY�	蛜������dd|��O �K�M�>�w��Su	��fs/i.:b�����m��d��69��o�',�io�?|�_8���'���g�I��eH@0V:�H$�J�K�!�� ��k�Kd�0ڊ��JS��8
�� ���	t�o��n���>�l��jl*g9�+�!MW&��Wta����>X����R]SG:xFL�^	R�@�2��"=�ql1	�JN�2�ƌk;v�Xu}��c�2DZ�@eRJ����^���n�2ֲ+���Y�m���R�%ܻ$��S�$��KM�r��2c�S80Sy�(p,E�@���w����d=R��ﾮT��]O�����@�p+d�i��nu2X�ݣ�{�z)�2�$|{:e��Z��__��{�R���<�r+J�U�۾��ֶ�NU��57YYf��J�W��d���!�"C�vw�%n��M�ju;����)o]2�{l��aV��bO<��=���z�6koaC,�D��ҫ;��D�:����Ǔ���c�]/KQ�8
�/���6�Xm�2LԒ֛�fCF�t�rtR�<MVjC2l�OZM�.�BQ��47���;-�5� ���^��luZ����DAm:K�P�Xn�r(�)S'ٶ�[lu���+*.P<�E��gE%�V���R7�X����o��g�-<N�z��9\J�x_�C�N��%^�Pz'Lc��̲Y�f��.ܖ��r�x~z�����и/��l*=��5���b��BЈJ|�?��a��qg*���o���2/��d�#(� ��Y�!>�|hY����(9�Hl#iq�U� Ƽ�<�I�>��N]g3',�a9ܤI-/���7�ρ<I��lҦ~��(Rat�=��!��|_P~A���;/?�A*���R�X�8��}AA�{�7�aK��z��?36����]7I��7�Х�^��@0b0���bvsɒ�}�,ˊ�Νg�M�!�:Lߍ���(�ıԮX߱#Ի�]U3�Ri��xH�(.ީSp����,�H�}ˋ�o���'�'o��w�{_�GF�8�&������F��� M��!�����/^c�RN��6ܵk�}����=�cǎvz`&�Y[V>���@�%Bh���a0�D:����?�$��G?���ܵ]x/���V+#��Y�F���0F3�����m���s|�����"9��q���æ�QGi�����d�]�S[k�᙮��җ���4�һz�O10��!�8�8���G����n�qt�g��D_�&<3������wD��	�M{D>C�����v�fb�}�Ӆ��2p�� � |K �R�~_*H�S4�1�X>�/^�|�b�Rƒ�g�Jx�����^X���mE�S�<M�͈SĻ�_|�?��O+� ��e�]6���B���&�������=��մ=�wo��cE��ED� [i?hA�C�� ^=�>r���"m�7Q���	�V�mΜ9�.]�t���௯����o��'~����a��團�[�X��J$�I�n̬�>l�u������X���� �"��%�7��n��q:}F��{t�:�,��6#������ҡ�Q�H�1��&�8���#!(��0�<������$4�&ݼCeo�l�s�;E�����km��+=�K5Ѷ��ؐ�l,^�:��z�~�!�/�"�8�d�T��X�:s"edIb()̽u�����]�� F��A�Җ�TY�V�c��x}����c�,c��2s�L:���[Q���A6u���5UN����3ֶ�R8�$p",#�1�L�V�Z���6L��(�Rٺl��}V�q�Y�뫮���fu�m�Տ;^	�=g�D�t�Q6b�Xk������f��*-Em�-�C��@ٿ�κ��,���
e$�u���fZJ��[���݇�zY�^D���zd8���؀f@�d�YnF������m������e#���+n�����li}�6!/�F����_~Ƕ�]jCd����9H��v����?܃���|�:�{���6�
�D~��g֕W^����CZ��d���q��ŀa9��p)��5��%\�d˘ZgϽ��s�|;����� ;ry�g}9�6#TW\q��7e�x;\
m��"���o]m��C�C=���~�6�%����OEn��y�w�A

ԕ��7Ѹ�?W%p|����C��< ��70�!�^0Ӷc�nkҕ��<��c>����3���81�̏롼�=ߢp����O�##FS{�g1��!�s�qx�ْ�;w�(�#����)�<b�``��a"�x(Rԛ�Q����%+_
q�D��;�&'��KhORHw�x�#U��>���쬳�t�Qg�g8����u#i�s,';�?������l���YL�1xgO�<(�����0������1�ہ��,���	c:��㾦��6n\�N P��Kf=����x����!��mCl{+��VU���z��,@����� #�p�A���'p3�
������ٕ!}��Fww�6����b�W���U�V��i3@�c���{�_~�hf�㲏�XҎW蒲�yx��N���LA�X��L�jvn�ꉧB�	�q�z��\��i�G؟���%K^�a!�th������s������|V��B��� �C��)��W�5�y�iXb�n�@�����&-��q���ݢ��d��z0�6l��|�6lZg3gN���F����[w���>�!���՗�)M����n����6�Fw�w�%/�`��n>|�E<]BK���E�\s�5vꩧXAa�dL��3%H�����Ó��qf�d��S?ҡ�H�����Z?n�=HK�.��ie��nQ�#��_2���#��{������1�j�û��=W��¼|#
r ���;h�nɸ�fv�h�<ȗ{�AU}��Gߩ�hqKKKr}}����>d��۷dɒy��s�U���
�H��$�D`h�����B�D�K�y���'x�o����u�\)C�{�c��U$�@����D�}��-����Nw���V���6I/������Ş@���|��p���������7�g	�����`JP2�B�V"92�3��/UX���K)3:�eF�`ԏM�x�#m�+���#GHydOF��]���/�g�^{��?A�B���N����3���G�G�ع�����ߩjz�߃�`���^�Hr�t)��� o�j�N=�N>�d{y�&[���Ɲ�+�:�6մ��wt���J,'#K�y���^_��W���	��|,M���uژ�)6��1����m}�yG���T�|r�~���Yy~�5ﭱ�˗Y�����(�[�Bza�eZJY�M�1�2��u�������d�-j�*u6u��ס���Ss-�p+=̲�ԡZ�����;����l�c�^�m���N�ΰ��2K++���B7�q'���.���ꪫ��F{��o�>im�BJ���V2n���<U�>Ϻ�S[��b$��Ofݵ�M�q���ly�e����^+-K�)F��Y}��u�H�T'[RZ�.�[���(.U;2C'EBJlZv��8�j�j�߶�jW=c�u{$�ԙ���Օv�aK�_z�.��r���L�(� {��*
^�a�pv

J�0�o�b{��V<<��3FէN�꼁S�b�������];�!��⊡�=-UF�NP%��h6�zu����M
)#�l��,�b���R2+�7���oV�R���s�@�������Q��e��Pމ�02�����=VT\dcF��Y9����֤o��K��b���R�d�k�����a���.�H�4e�/�x�J7��O���3��P�x�w!�a ����6bF\.��nUf<j�Ȑa栵Âը�PSF%)#�c��k|��˒=f�}O�d'8 G��T��J�b�����`�z�TF�}FT4�RI�1S�~7x��ϝ;W��4{��gdo�sܘ9�ַ��.�o���4�Y7���R��Fh�8�=�� ~Q���\���6n�d�$�1����W^u�e�͗+��A)?(��5��	��r(fKQFI�}(��G��8����	��<C>���xN�e�`t]B�}ɳ�eT��
�m����p��>���Ϭ`��g�N�/)��'� *��
����#�����0Q܅�~cLS�8xIPU\F�]�4`�����Gx��~�� c@��l!�x��AI�\<��L�7�����~0�tP�)'���NY����rc�K����93�@���� 3J�^v��޹6�g�'z�v�t@�[�hr�w�w�M����{��w
Y�`�X� �x�> ܗ?��C����Vf8)�8�5(����)u�@b{��a�4q�0P\�c ��
�{���H�1ڋ��n)�fh�;e�/��
�0H�>,����B%C�|`o��^����JY��D�g�B}V�ڷA���T�ɲ~=)�g��e���OBnC��p�H��?y������.�C���/����r^F}����H��VlS �/StH��g��Sf˃��+Vl��~�7��������S���
��S����_���˗'�7��p�NX�
A��>�@���w��|j]���$��	�������9��ر�8?����Jʊ���SG?�GQV�Z�ތ�8�g-(��$�#`��&���p�7���@�������@j�cN�kǞ��^Y����l���~��<۶V7�g6�֛�n)��+{�z$(�,Uy�ґ� ��n I`J�Yِ|;lR���d��l>��?-K�C��C)g=��o�$<s�T�(���Z�0&�7�S���$ː�b[Kg�ʐ��\T %2Ye���:1��i2�T��F��U�6kil�Q##"?��ڲ-��_Ϫ-+7�r�3�C�ݣv������:�Ռ�T�d���aMR滛��W�@f��(ʔ����e-M�N�D��/ET�[C�:&)/�gr��(�3GZ����Ti�f����[����m����k�O�aW`[wl�$u#Jʭ�!�Mr�[j��Vfի��e���2�6[~�t���ӡT٥�.�_�
F�����E�ؖ͛]��r@�
��v�
�G��?0�PH3��5bf�4�64n�x�A�8�$JRlÆ5v����/�,%~�{۳��7	���s�P�0�����M;��E�8-���e��{V��ک:�}��A�`����b��I���)�:ƏgC+�� bVd��Hs蠨�w"�}�gt����g:��x�͍/]�e88C�g��	�0����s���Z���@Bf��0+�c
f�P	���X��R^~�1���$� @���
FQQ�B�w�l�F桼�(�^�� ���QG��0�i����&��A=?�S�Jo�x��h��R⮷�^{�O�gO���o�<�{��a c���.t�dI&#��lQ��*���?�r�"�%�����}���w���#�8A�������S���rEhO�o0f�Ԡ8D@&F���i��
�~���%�I�Ay�����&q�*�%]��7��to��Ӯ6h_3���.��g�����2@������{��� 4G�(#� �#��W�����p��Wh��~��3�vS���{k�=} Ye�.䋑�%�=]������	M����� �7�%��B��C��� ϣl�/++�w�~9���b��`Q~���Oxm^;�@ucI8������ �J�A��r����~#��/]�T탻��f��G �e�e �Ϯ��]�͐�D�{��8a���P<���
�Z�^#^".���=me�+��'������U�I�H�gZ9=` ��q���0���qٛJ��3x�6�C:A駞ْia��q���["����@� ��uh��1�<� ���:��Q
�ƴ�&QN�o��y	 @��d�y��r�ʍ7�p�u_���_�	�F��m��(S8���U�V��_U%&��'���� ����aL�EYc�*��4>�/(ҁ���%��e��j;�ow��w(��r����|�iS����/�`�5�V(%�E(%9��P����{W�PT��$�G�u�J	UaÆ�]��V��mS����bkh�P/��P��Kኍ�¥p��p0��]���j�jhy��W����h/?�B8l�܂b+���R���.)R*�����Vk�oq��戱K�pH�e��Z�:���TkS�ݯW��%6>�ܬW�LF^����X�:�t)d)=��ٮrKq�J���.�O
<mZ��j�E�YZ`9#�-)7�d�X�e�h,J4�F�À��\��ɶ)��%�VV1�JG���Mm�)�Wec�<Y`���K�L)���ܥ´$+J벉���Cw�=���=��I{��g����N8n����ڷ��O��yK
���S9҄oa�G�+��Vm�m/?e�m��'{亝�N�b_���C19-�N��ԡ3�"�,D�	/D~@!���rΝ�},��8�`YKY��!�(7,?�"#��������KKd(m�<?�Oڱ���`/���Ǎ7���/x��I�̊�7�+�;�2c�R ��ٙ�Y �.<;(���Y�uV:1N�������d�3�Ɍ1F^�X��{CT>8*+��6��Z�#� ^B,G"��z(��JY������3dMh�Ύ}A��6!�hkh�o�G� �P�⡪=jwʈ�@W�$�P���ߴ��ʉ��cf�%dٹ,�p\������.�	��]�P^F���>��:����V�ڝn8�u��e2����g�����;F7K?�F�r���A��!�����;��������o�?�]��� sZ����D��o�Ӿ����c�S�	���9�r%P~G��t}ҿ�3��|��*�a���~2F���@���j�O�z���>R�%�8W�$�'`�}X�����;��6�7m��=���l�<�s�>��^9��<�`wj��Z�}���g� i18IZx&���<)�"fP�G��yη�����q��A���2�r�e��(m��\� ��?��{����L4/��!3}��q��;8h�� ����|��y�n��s��o}�^|�Y��4;�s�¾gx�	eg���y欙~��gBq�>��0��_�vw�!� ��'h0Q>1p . ��n�!z/QFA���=8e�7����y���=x����m��^?�VW'-a�,e��"/�$�������f g�}�o���C|N�خ�����{���b������y����q�������,y��j�6�]`���i����\u���~��C O:�4;񤓼�d��"��
@ ! tz,�����!���(ӦN��Yb���k������"�#bB����?i��V1}pƲe�V�H��u|9B�%��e���H����o��`���#������D����l�h����c��-ߴ׶����\`Y�����_��(�>	��u`�)C �O���Ce�B��W���'����&�Za����Jmܔ)V1b��vX�:��:�dkR �]O_�����E��(�,�h3KS瞄��^u�2.�o[s���3�0ȼ�~�L�,)x�˒!��^oeY�6e�P�ߜd/��e��f�)鶽���3󭵽ߚ�p� �GB\m��T�����d�w�˺��`6-��:U���&��m�,�>3)]�f�K��&7YJz���[��R��M�\�Ɔ�tڲ��hei6j�T[�f�m�i����نO;Җm�k{ڬ`�p��ʕԗ��E	zJY6f����b[y�O-�n����ʀ�V{l���v��g���{更'�xڮ��Jw�2R�*��qD�;Zh�{:(:V���ٽK���3jO�Ų��,*S��KB)�����M�O���Qw��%Ky.+�Ǡ[�x�~�����Ű|���lF�����<�b�����0ru�#�l���w<��0|;M�>���3�pG��kT�0
�h%#o�	�FW_�#:rff��{$�F|P��0*��F��y��*U������Gi�5��j"RFrQVb:ٸ�L���'=ڞ{�!�ap�=2�bӦM񶯯�e��uKd	2�M9���E^,;��ϱ��n��>_�2ă'�8����`m�3H�F7?q����f��������=s8���3Cy�]�@]�]�,�y�;�!��&B[[�/eb�	C�B�B��ăeZhO<#}}ʌ�F��OUe�-^��}�k_u�-�9�p�#|'���� �g�9i&>��O���Y���q�hV-�PR>����Y�g���Ӊ�H;�:�;�^��۶��������j��bx-O�v�c0��=b�dxҡ���3�#��y�u$~��y�G#�`Z�'J_��Tx���{:U�&wG~�ɧ�Yg����ۏ~�c��(�2������b9�wl�����Va?������^��9y��̶"�e+���'>�B��)��3�g�0�2�r�`g��=����Ѓڶ��-S<�<&�?4ey"���8Ѩ���K|�^8`�9�3}d��ʗ��- L��2����8[����w���N����E��'��!;h�8�!�Y =R~�(��z`�Ѿ� ڂ�i�B{��H���� �~l������B`�@��ǇpClop�5�	<�wB�pe7ߒ�#l߃3���2?'[����ڵk��Czח����z �>5�n�s�Ό%K�,�|�;��Α�O?�ē�.�N��g�u&��ccjrS`�H�HqDb��"��&:��O:ŉq��uk�!�h��Ɔz��k��}����!�C��UR/��b۹c��3Z��qP���&?��<c�#�r�w�C��
�2��\e I�ig�	G������[���#�
�oɹ��٫��8�\��v�0��v)���%�Қ��f:��n}�k�b�VRd�2�2�r,K���b�U.����Zd�I��$[������nC��r�2�Ġ)��I��#����}z���v�/ȰaC�0;Ͳ��u����QY�k�lX��5�������fOȶ!��xy����YgG��l�f��v�x����	_�/5Y�'�7��Ig�Iɱ��,�[Jf_�%u��2����-֛֥�'�&V�[rm��}�Qkܹ�2:�ٸ�t��n��sf�ʵ�l��7�֪;��K-k���)�M�g,��B���� s@��L��#ʭz島�_Yv�V�m���.W�X��G�{���w���=bW��*�Uff}��Hw�?W"�;*�Y�͜a��Gw���I��+ދH���H��*3���A� �����}4Qq)O��D�!#�	<���D<$F�)'�%�+��/Fo"���F��G0��>�*58�˧|���`���ع��t�z�R6�/~aϑጦ�)�`��5�'M�2���4~So���1������r�&O�=H[�l��GI����+�*/�D��K�7�ߢ��q�b�1z7V�u�;)�]�_��B�-BQQg���Sm���h������9o)8E8h Q���/��Q{G�	A���`��-v�ݿ�o|�/��C��g��[�9s��k�yO��&E��Q��˗�?Ս�l)�$�$��v��e�q���Zu����f[�l�m��I�g�H�NW�T��� �$@�@�	��S:��u4�#�1��qX����	�/C��&N�hx�d5�ZQ���=�kV���S�s�7��V�m�+Ȋ�LN�O�J��OC�( n���N�*yD^��@"��w �r�;��۾�nWb{��,�&��`;�۷ˍ�?�{�s�Q������~�S=v��
�?� ޔ���]�[�0������~��Q��eH3�Ǻr��.I�fp�L����d?W�}�=f�/	e�8��t���΀�/�U�zhx����6?:����;�J�����2p�e�7!���~��N�t_}u�珻���,��e���_�&@�#��7�d�@(+��Y ��83X6\�ԯ<YB�!�l4���6���K?��+�ӝ�x����q�$x��	��1���46Hh�D<�s"��@�u$�؆��ئ�� x�tJ;h7��v#.8$���F���=�m�w�w$�]�I~��[����?�����[�l�Rx��鋷�~�lF!O���9?xva�����#Q��Y	H��H��	��HX���?n��uϞݮ((����l��q�|�;/��n�O;j�����~`&^c���4q$��@�\�O�X�X' )�3��F�����Gl]�-v֙'��#��s˷Z�Z��c,9��:�$�%�3d�uI�i׷�Bܰ�(��QT<qO�. ӳd$��m�:�$1k���VXVb}i�V�:�	�%��lOu��n���<7 �p�-��������j)���L
$��\A���:*�
KS��Ɲ�����m{�z��#MZ����JR��ն�[S{�;{�+ʲ�����<ݗZW��!aߪ��^���ӗ���VdH�����g��zSWC�ijJ���ذ�t++ȳں.۴��z��l�!ֵ��|�+�i���e��=g�ˋ쿾����SS]o�^�Q{��M�9z����ІN�e��)֪2��	ӕW����#<#զLc����g~��k�c��R|e �����O?�$��G�����]*�@��(�؎�A@B��<u��-�^�-�"8q�,�����>:M<6yBq(/t�.���M6�+O��#��.�*����{�E9�����4���!�9'H1�2�AW��}(Lr ��q�]�98z���e,�:�f�/�Ү6D�A��ț+� p�o��q(w�6(;J��t�Np�;z�H�3>��F�X�ʷģ\�e�=|;��M�*��|��Y��oݺ�֯_+���T=�;�#���ߊ��)S����$���{�57�2!"�3+�!���p-~�<���P�����}�k���l���~�1gf��#�6��u�[�-��)=z�~�G9�+"^��i�}�'@��N@�,'c�:���=�)��a�e��$�}Ш
������Aω@>o���(��D[��|~9H7[u+����ϰ��>��1��<��~,�o o�pnJ��y�\��.ǟ|�	7F9ӌ���|^C�p�^H�a�G����ԁ���H�ĉ�&^b�y�3�K��H������R�p���[m���_��n)�\�v�}�S����,����By�qL2��yy���,G���P��O�p���g����o��A9e@ �f:�ԇ��T������lJEy���K�'.o�O(�>����8ԛۈz ��1�`��g�n3gδ%�ݦM[d�!�H�f�A/�e��@B����G��vD��}��%Ί3����C��>�ʠ
��<@�|�á��bo�M�1��ġ޽����aĕ������W�ê�zz#�����C��/o��H� ��-�3� �i7x\�|���廈K�!��!W�A����딮R�ν�����?��O����(�ކ���?�VYY9^��˲-��5]�n������HT�t����'(S�ND<�Ӂ@x��� �!e	���^��6��v��iS�Or�w n���߹�a43�qtpz<�DH,�����%������$�ۅ��y�:QF��cÆ��-��&�f��2�M������/�R0�˲�p����=!��O�.��Ȇ�a������:�=���u[���NM��,���Lσ����uq����)��kE�}VQ�l��شI2��ut�ڮM��:[�b�m�^o���X}c��6v[R��Z�vmu�U�uۖ�[�~���j�m�j�	��V�RJS~Q��e��[7��Ԇ�)j[��{z��\�b�����dc����y�6zD���_o��-;��F����'���/��SG��qC��~�;{�io������mŚV2b��~R�l��	2^i	-��+��]���R����ږ����*+,�!��Fmni��ӧڥ�^�4pJ��W�I���G"�D>�4�%�� '\�"T��a9��y����ٶ-(�a�����]��=K�2�92�*�Y��� ͆2�w��L��cP����E�1��ϡ�!݃
jjv3x��^�H[�P[���C1@�F���PxH��aQ֠X#N�� ��Pf��'�M�q�������'	MM��7�� �^*L�g4Y���QXf8���)�銗��Fkf>�>h���� #9I�x�7�33C�	��G+���Y3�΍N�� ѱN��B�Q���~�QG���|�5����	m�l��G��l�ƍmÆ��m�V�;q�7����Ey	̘d�#ݗB�!Y��a�.���T��l�˩:��%��P��7k7�o����{d?W�����}�{U�;��s��o�|�v�%�l���j�\�?�6!/�+�jϞ]��Ro�RfH����Qf�Ar�kcn^��YaG=ߎ?~�-8j����7;{��?�|([��J�'�C(����lhl��ksޡ��+�G��6��=}i�a�#�48IA�,}�����_��~��˰�!:���3��j�Ӏ�܃-j�Ao�/�~CH���V�!x�$���u���D9�3��I�3��M��C޹��Yu,5���0���@����D��/�=���+,�͛7���{II���o>�-��ԇ4�٠����e`ڃ�h+"_�o�Ϩ�v�.����>e�1����l��,�mhl���*�ybЂ�ɬ^ɊNɄ��;w���~RcY�5����Bb�����"�ߴ�b�x��ў�7t�s���Q���`��o뺺��c�9澧�~��=H�� ��x���O}��G=|�-���/�!�r�0����y(`���qsC4��΃��! �H$>�"��b�����$A�V�?�H{׻���;�D������嗿�G9�Ep���|c �CC(�AH|��_2���/�M��@�@�Ajo�3O9���[`O��f�}��?��(a�}b�	�T���¬Z���LON~���}���Q/�K�Bԯz�}m��>R�q�:���2�mﴌ�2˕"���i�z7n�:�HY����j�-R,��Y���^��'%&�J��� +�r�R|�m��]�m�.��i���l��K���|��	�L��i��2D��4�ت{lۦ]�e�f��LKΗ�ԗj��Ce��HQI��lfDy)V]�b����BJ�I�'��V�W�����ءy6,[�mk��\���J��-g�i)��w�`���ڵW�kŅ)�n�2[��5+�ϴi�ǻS���o{Z����d��n�Ͼ���W�KQ�d5�C�6K��ټ9ӭa�{�;����m6rg�(����s؃t��5����.�ԗ��p��B1�W��A�%?�$a����@t�'��羧N��g�`S4 Z�;�8DE���2�,�Aɪ�~ǼyO�Ĳ��~ϻx�������S/C�~�?Sڑ��O�"$Ӣ}���(��9G	���(霵�b��I����2�
#kZE�Ȇ�P�1_���W	���]�<�! �3Si�� �)�5�G��%���E�1r8�j��>�N�kk�}=Ȧ�#�B�3��V��`���e*�V�40LX
�cԐA ꄬ$O v���׿̜L߯Ìg���:��c�+8Ha���<C�,{ n��?��������W\鳝,�{���=��'ҍx����r�vd�Y;����t��b��ˠ�:�Ccr;��4�0��!]��<q���� �O(7�V�8!α��}N9�"�;�R�����Gl�uk�Y{W�;܉�cAA�M�4�q9dHXf�`u
!��e��}�~��?ڣ�-V�z|�%�N�QN�e��Zѯ���=\�ܻ��s4�qOna暶 D �$�]$�N�
o�GcЉ6��9K_SR2l�(�le���<�B���@[C�B��s�\0�~Рb�U"��@?qXt��Ez�{��������s�4���'�O�[�B�!�~��"�q% �i������*�%��?��h�Ƚ"����{��t��%�J̪CO�frX�-��=�ʡ�!��<�$�@�Q&�e�;aJ��*A&ц�e�]�W襦�����{��Q����v�O���>�n�l+ر}���6������̔=�0�����5�f�����q�<�m�s���7����ox�g�:��T�͕86�`h���O|���ۿ���� [�߆ȚM���θ�;��cJ9��k�E,!
F��-#8jx�
�e07�(X]]�'��G� @8��Ie�����X�L���c��3O�47o٨|��SO���L�Ӄ��W�G½#HR�N��	��{uI���I�)I��/U
_w��u��i'.��ga�l�o��,�b��f�X���d)tiRhṤ�tXJ[�e��Z�r�R�դνU�_uA}��$�n)�fȨ����g[�n���VY�p�VTb��G[����V+Yd��b]�V_+��K��tZNr�1<�ʆ�X����;km���VW]k�M�2������&c�2�
��l\E�+H�ގ^ki谁�d�kl��$��:rlϮ���bU*cM���"+.�J� ��d���(�Ԭ��벎f!��K�rj�e����(�\յe{�-j��_�\i��Ӧ��η��f���-�z�]��VR�a=�5�5ڥ�m���^[mO-Yi������q3��s/���~�6M�c`�T���bS'���+���Ko�e��0��5��L����<��3>��$�Z�N"����-���?�;���C�+����F��o��gF�V
�14iވ4�t+z�?)$�FQ�1*b��~� ����h ��@"Y�
ߒ���@�@�1�b9�}bP��ㄎ���(�Ç�����H@����#�V������7XN����_:�'��A��%_/�`9�!�7�+�ÈBz�,3I���1�RSS�\�#ڒ�X�:>�����[?gKJ..Ùya����S�Ѡ�XN	�0"�i�t���h;w챺Z�Oϲ�\hR��!:l�1��@b&��r���>v�}�K_r�:�-�z1����"Ƿ��1�y�x,���s���������Y|K Glϓ��9o��ּ�� oԃt��EU�D�q�����ƽ�wy������%Ə�{�����e�^��򈌘��@�𧲃�hF��"<*�	x���G�kW^�.;��|�HԤ��	{
��j����������tP&�"��q��bL�X��@+'X^�'W��v��PtYnF`�����S�.2���+<h��������Ya�������bu������JR���
O������A9��A�s���1.�fR|�ۃ���M�'}2�I3|C{P���2��\�mJ�L�^���=���.~���=�F���yw�e��QGe�/�6:]�����wk�0�]�i�N�3<�L��&OT|<�rVd(�p�@o��\^�Bf�Ox.��c�%Ǎ��?ܷ@˱�uu��&M��͊������K���ʹ)^���U���'���/~����1�z�-���o�ئ@h��"MqO��w��x�v�'��o�=�g�7�D����s�����N�Fj��m۾䓟��n��e�@�m5�a��0������_��W>���׎�uj�Z�5�t�4��D����NJ��-�xfu��0Rò��#�r�{���s�CK�]|�Evʩ'��n�*9�����������o��`��A��mȇ4)*
�/߃�)|�VW����@�1�����(0�'�5,�ڤ(%I�>��l���-5֜^n�#�XOV�u�ANhF��8��O8S��� Mƒ+&�f���{_�����}��*�g	��R"7���u��[za�����|Z-)+�&N=܆�Z^�:�����#E5��ʇ����V��c[�햒�Ӳ���ȩ�m��r;f�DU�i[��S�ݶ�蹖�!�O�`T�ڍ�b�Z۽�JFa��=��{�<k�_��Ҷ��ڡ��m�j�s�Km�e��H���8tH�e�XcM���5Yq���������}e��{n�5�P�ͭ�o�(���a�G���~��ַw�]ɱ���h��v����w��;��5tg��~;���l�q�ێ�&��aB?,�g�;����[Zbu˟���e{�Za����k�^;����w�����{�I���K���@��)4m�5>�q\O�8Ѿ���JA�k���/졇�)S��� 1��A��,~������"=�%%9J3/�����HE)���m6n�9�97'����{F�鴣@��TF�P����RG[�⑶�f�s�,��#��H�h �Α7 q��	#���h���R.QX�1�����C���8�%d�3Im��TgO�F�a�?|JGDG���L��,A���P��>���Uo�1jϲW��a� q�ߴ_�r1�E�PJ('��yF��VE��x�C�0����B��̜I��!K%YE{�3�e'嫭�U���d��,2WtU.?lP�;���b����^��w����o����G6l��܋?�a� � l�l���?j(����V�q03D�Ĭ
 K���]f���W�� P'p���~� W�1�.���XC��&	�]R>p2�,$��t!��k�7��Ni�>2�.�7��yϵ�.��}2�������Q�lq�SVV0��v����R8�/����l�om6z;��qO���:�N8q�/�qM������a+W-��:�6oZk��G�_�퓖#��=vjZW����o�}z.����) m�=�^�j���۶m�=��I�=��2�I�}��>�>s�\�}��������v�5m��N�W~�6��z\��}��"V=�>�;�,|C"���p�0�y�2�]��4xC�Sb >���^w���h���{m��u��9
=�e�ȟ�EV���U��d����<$_��q23����kȇ���_(+����]��+St�+ޡ8���d�e%^SS��ر�^�����'&N����spZd6m�:�|��7m�p��Ŭ�!��;������_��ӗ������'Ю�f��x��,���V�Ũ�2�%�y�0̽����+8�@�!c�a�>X��U���[�>!��c7�t�F�� o4K߆��p��7��/^�j�eee9t�]R�Z,W��=c��ϕFF�\���L	�m��	�N>��1Rƨ�4������[��E7�N8�s��z���u�w�^6O��*p���p���8Q��׿ 3�_��pS'O��#�ض���J���m =�zD�$ɀڀB��q���Qz��_�Q�H��i��Xg,��o���4]xj�Q�^'Š���/=S
�����7���N�׳^{}���u[l�����b�F�y'̱��9ܦ-��tu�5�a�2�L��S&H�֫m;�YJю[��VZ���m���Ͱ�ÇX�@�{��6a�M;�pϽ�v��L�ge�tw�_���R�kCJ�mXy���@jm�-��kϿf��+L��,����G���,-,�}�vX펍��s��~+-)����}6j�Xw�:y�t�S�nO.~��G�Q�^l]IVY����
�¨��P���["���Vo]u{��q�X6�r�g��ߎ�E�\���߰�~/�Ze)\����F@��+�t��`���駟2���YN��I¬��M�fϔb�����N>�4��۬N�4�&Uf�y��)6�Ý�࿰d,x��;��oǁ�m���NOh<�#�?5�o�P�A{�@�&c�r�I���:�D?z�h+-+��^%���FP�'�+��G̜�D����<A��=�Q�G�A�8Aޔ��p�cҭ�c��<3H����V���+6�ӱ����1��-�E�PD��B�cY�F��=�#�5I�Γx�ԑ�A1O�E�J��`|P�,��X�ܕ)p�+�DF��< y��S��L�����Ou���0��3��Q�@3#��T]�=M�!�\�ڽ�q~�5��>�A;r�|W ؓ�$���iӧ����?N�$ۙg��1y��O_�&M��cG�?Үz�U��U�WY��P$�0��N�j�jo;�:��M�؞>k��W�f�V������&���կ~i���g�����q�<��(fe�5��1sƊΣJ���V:��O�Q��N?Ѯ��j[�b���G?���^��T�x.�1e(��zԶn�&���=wW_�n;�؅q������Ea���ΗLF�!�� �>��l8�`kx�2�O2�>8tK>9�y�Q���N���:Ɩ���mܴ��`H���+qV:���E�@w��&�97���`�ȃk�/���m̟�9�nx�7��;1
��OL� ���'��� ����;w�M�4�֯�`���s����=F�@�B�<#@gQ^��M��'|�ù	�^����}�L����+���f�}��lmٍܸd~3���[-Z�;ɵ��!p�eW���gw\���<��� ��b�4�����H�x'O��
�*1�>'��]0�C����r���r���?*B�uD��4 ��E2�Ir�Eߴ��׉G�Ԇ,U�S���Ҫ&���Dd����A�wH�$��d����ݓ.|����Y� oH�dp�e�,^����۷O��	�ĩm���D� �@"���!4>#.���(l��'A� �G��$�D�q]�[�֎�;G�Y��e�3_H;Hb�3S��� ��_؄:( �s�B>�{y"��AH�����Ҵ)��b�(۰k�5t%Y��ä����#o���݈�S�Il�A	x gJ�[�q�3	@�KsF���+.�v)b�{e\tt[NQ���tkm�a��dS'�ZI~��X_eK�UY���!�=v��#mщs���R���l߶u�g�k�����>u?lx�ѵ�x�B��U=d<��J �Y��R�H��V�~M=-���b#��Ȉ�0�pKKN��M��)�(����ѹ6mR��6[��۰v����d"��Jh�c�cGY��s���q�mV-�ߧ��E��i��,,�����}��f����f�~���:˶�f	�T�m��7�̩8���cyRRzj���/Xk����@�����F)�c��K/=` �Z��$�DJ4�Q� @�0�qh>n�E��9���r��Q\�!08m�t�0q�h��;	��,�ݤ�b3fL��G)��=1g��b�A�ݻK|���i�����^7P�݀aC��7�(p��7$	�&��D��m�p�$�۱���N�F��d$t���^6�3pB|�b܌��D��6�әG宜�(|�뛳���I�4�Q�ǱL ﹏J�cxS��2�|�GZ���hԠ,�74��áՔ��)'t�K�ŋ�0 ���&��(�� ��Qe6JG<0kF(�^v�L�h��l(��js��v������jYD:G�� ��	ޮ/����Rb�b��S�EY�-��5�����B.���t͵���oG��N<�x)�l��c�7�`��p����駟j�k����=W�Yg���'���W^y��{��v�E���	'oG-X`�/]�4Jۃ?����)S����c��f@S&�'q�Sf�z%-z����!��&��7�n���|9T~~�/o�>}��/{?01�0�	,���Q��˘���G�a	���w]y��|�G�z����k~�ēO>m�����?�Ǝ���bV���P��|��sn�՜ٳ�tB-���w�!C�W�裏�ku��1p��gx!�W8H�/���/���ʕ��i^~dM"~"� \S��8�x������N�N�,Ńv �|�����<���,�@e�b ����'h�2^#�X&�I,�A����в���Oi1nL#1�Ā� �'O�t��$�	ƨav���2�A��}�Oë�j�I���A�}�C��!�y�w��@Bp٧v �<'N�dK{��'-d��y�%�\r�w����:�������x�g�&���$�rR�X�C��� p伬+8�k�q�oc�	��押�8gIt��Y�<�ݻ����wߔ��_�={֣#F�xUx\&����3g<|��y���YP��=t���Ξ���ֶ^�=��.�g��N��N�M��3++c���f̘��\����o����m �������K���iӦ�j�t��u�a��A!��� �RD��'@PhJ�����O�3����2>�b�%b����5�zl7��9sf�3\�[�f���O��QJ�R�F�**G�P^ʅP�>;x����)i<�@JV�2EJDiy�m�[c=��V2�0�Kɰ� D@��~���‰σg�I�ɬ�P9X��#�GP��&�H]��#�X�]P��Lu������V�ξMZ�nJm�u2"�0`����򕛭���&�g�E��9GN���6�߾��m]o=�Ֆ�I[�[Ss��f�(��O�0їS���U�`C}�+{Ǐ��#�[[S�uK�n���T�߬��*J
m|���Js%�9ش����^ f+emڴݚ�[Lv�@8��W6q���6UB,ǺeX%	o��Eơ�{�o�=�XFz�M��R������������_�Ɇ�9�f�x��ij��]q ����R�]٩`)���/=a)]5VZV�m�gA��O�Ҧ��="[�n�{�x��a6((�a�>��e�و�U�(���sf�M=̕�G}�V�Z�V̎����M��R̷l�)^0�;w�+1]���)�������c����Z�\B��0���p�(�'O��B�w�%�\A���q�aӤ�f���*�MZ:�s鴥0��_�3M&#� �#Pox�zF�.���TysG��G�QD��w��x	�2#�	�����
��DI 0<Q :��/��E$��r'�޸�H:�m��^x�Y/F�Y�o��rbQ7� P��YGG�Y�ΰ\���Xp����T��e&���E���y���L
���ma�f�U���ԃj`�R����A
�8C�ec��WF�1��出R/�ĳN8�ޱh����w�a���x�����p[��.���d�3���L��Γb�����=R��o�?e��􌥌�K{��[�H�;ҀN�,k�]t�~������W{V��:9·�A\p����w_���e�]�΀.�x��iy�P�C�V(�v�׫�)��c�J�juzmmk���j�����穟:�����~�֯_�=���],����f�{f�0R�x��[����;�N���z�e�9��'�#������L0���^���8�Lo����U�<��{S�H
�x�{UVV6���?��a�[��D\G��_���τ.f���/�g�a����5�O��Ѵ+i�o��ȗ�7��ybx3�e������.1�;�ź���y%��Y��X��ח�������qF=�4��M����K.�oU��H+�E|��op���%�i��A��IL���mY�h�����¦�C����[��C����=z�V(74G^������o�/����֢l�%pj�~ðG��&�+c�a޼#�Ϛ9����>�K���g�q�#'�p³�/����;wΦ�/ǲѣ�Tgd�%�8|�����V[Wױe��d���Ϩ5jĪ��������c��qK�?6q��G��/����$����7@hѷ���暂�^{�7N���t�8ୈ�t��`R�M~�����0���P48����%K^�QD�ą�*(V�6or,��N=�4�Aھc��FP�a�v�7�:��T9 $����q4��<0bν����I�5������x,�afd����2�U�b�%�=t�u[�u��{�%˺��aI)2��;%O]����֣��"K=�14������w�)�w���6�2U�����s
��|)em�u�vk������S���3�[j�۳~��W�Q!:���ѡ2����E��G�6n��^���zm�����.?_�=RSU�t�M�p���bmM��#� �F+�Q\�t'�8�-�klO}����ZG[��wvYj~��0j�x�S�w6�ZZ�:�.)�9�6�b�e]m=��3��sϾd����^�����M�{�-<���~����R�Mj�8�p�YM˙+I����"Km��-�>m��6c�og_��0k�lW�2D�@��,�/�\��mō��+�K����8J�	(�t�z�b�J7�|OYV���Pjc�������v۾s��T1r�������3�;׼yl���~�x���"_B��v�-�ا?�)�]"�i�믿��u�eR�����>�n��7�{�y�̕�jB'�.�;�������s�*��8��0f��B\:x��Md��H����[f<0,�7��Æg~Sǘo��Af�A^?�,�@\�Rpx+y�f�j�ݪ�+el�(��P�YE�Ӟ��Yf���� _о��\8� A�Q�u���N�+�MfOq�� =�,p�;b�
:��k����Z��u���r�_f11ή��z(�(�W^y��3�(J��GiC����$�?�����%s�gmf�P��F3����+�d�6�7L}�%�ꫯ�L����|֊����z�g9^^�=��c��3��5x���z�A8u<+ �6�� �����5�t \�D������iӦ�;f/��N��Zᕀ�~���7Q�hgރ_�-+-�|���6䨽(��!C��$_Z�l�
�S��'6o�(<�˰϶+��ɓ�yޤ��Oۊ˝&

��]W��&�O���-[��[?fw��gN�ű���i�K/�\�0V�H��@�P�#F��óɓ���4�Ҷ�۷�� ��SO=ew�u���t|s`0K ���sϽ����mB��q��&�[O�<�aO]c}�ʾо�����=��>��22m��5�7�,�y�k�C���B,O�?\i��J��1�C˟�����	Q~p���F �g��YOw`�a9����@�I�)��U�FZ�� �@z�L<��r}F�A%��J�%Ҝ5���W�J��"���^�=[.�dу2��I�P���ה�w��g*�	�R.h"�|�@>1�����̀��zL�e�c��%rr�ۏ�7����G6��4�?��S�����)���ǣ�^�d��{����}�{������u�u7�nܸ���� c�����{��ƫݳ��؞/�#�e��&�544VΜy�/nzߍ+�|bq��?���'��{���~򓟄N�M P���O0����-�� ���	9P�H����A<G1����_���1*�3��t<M��[�%Atd �]Цb�%�%/|��@X �+��\
 Ba��c?OaА#�p�N���p�C��t�?���s~M�x���n� #���
UW�%��D��F&�����Ђ�S�_��!�/#Kb�z�M����2��*&����m�)��Ql��9���m�'��;�S[2`�_�]�VJ�hW��!!��^�"�+*/-��}�����7��5�u⿸��_Y��q46��6W��T����r�Vjj�e��J����Jh�g��:�1E6�(�r��ު\/� ɈL�-����1�FL9̊dHt�tXS�~�ײ�Х�U�5ZmG�M�j'�p�������잗���.;��s���/�Δ�M�'#�����P4�i,�huX��|��I�=2�pE����n=�@��: ��5<���+��N3*�����~-RV�l������S��Y�\&���OR�mں�~����?-�:}��3V,_c�ʰA��n� y0C���c�6����0� 6�Ǝc��G�UO��*7������@>�+�j���.B$y�Y6�r.f���A�C�|Eyǳ�bX0G1�{!<���q�" �	Ȯ(�"D��z�g�D�G�g�[d�P�@;3�����k��ж���Z �p��2������ev<'���=�ĕ8y�eb?��@�݊�,!�W�e
��9���3ϔ4�N8�7|pq�Q��A�N��Q�~���z��+�t������G}�~���ؗ��ew�~�{��������~���w�B��˶v�z����3���=��f�k���"�mf��N#�e��iOڎ6@SG~���6��@����3�K�|�Qp�LF�G��{mm���?�޻���|�=��#�t�����y�)v͵WZِb������
��1��n[6o���L��S�l����܄�OTF�gXE��[sÄ��~ĩ��׮]k��ηd�-UL<NrnG�euǠA{?�����iF��w������'����p�J "��/x�c`�.�K/�T�yX^`|�t�Mn�1EC&�������*/�\1��@�00���c��<ȀH�{ 1 �ݡ@���7!��6�ޒƠMXҋ���^�Z����`�g�́�q>�Fc.>C����=m,Ň��f���1 ��3I��e}TZ�J޽}�)��n�0��& �L�(`���(?C��<��!��,���VӠ�Q������o�6PW[S7}�����z�>����s��'��r���MMO�#�5;��q������?�}�Mx�O���/�駟X�����~U����0;;+G�TΦM3�y橾����I5���b4�~�**?1�;>�}$�77(�(|��=tXl� 07��{���	)tp7](f8m�e���W>��1��*[��s:��#ƪ��lv���Yi� o�$D�z�F0E%�4##�B�12D���k/���E%!����O���X��g�T^��O�z7���N���tI!�W_m)9�vؑm�a�,�8�z:j-����ȳ�Ϝo3+R�a�2�ٱ�z�1L���@H�b�B�p�ᡦ�f���K}��R��T��L��~u�}��t�Ї�j�p-�(=c���0���4XK�+Ij��Ǘ�Ēt��o���d�HSR,�t���>��G�Q��� �T��Yi֦~�O��V-�f�:�ͭ-V<g��tÇ���QG�n�cg��mնv{�{	LS�W���
��}V���^����57�ۊ�+]Q�#|,������F�7h)�h��36 (�N�99�i#�[���v��,O�Yp�Nz�W�5����Uh]�y3��,Hlō,Fs�����|�Y�|P@Y	����ڟy=��hhj���/���/iBQ�|,�do�ţ�j�^꡺�,1��� �ǎ�ߑ�A\���B��ό7�G����0��l�u�`LzQ�g7����V�2&��&!���58CiaY��Gq�/�#t@�(;�.t��+8��H�tH�o��%\�7!<�M��{���RN\�H������j��Y�ɡ;%�3S�4ȋ�E9fv�Qofw��%�co]����쮻~-#��2z~�ׇz��~�ou��W����z����?��=��Ӷe�v��W$���Q6q�++f�9��1ߎZp��#L�X�Ø�B�"R?w��z�s�;���
	�~ 0"Q6�'�|�I�q��yGXYy��N���\WtH;v��3e��3�-;7�ʇ����� =�N>�D߃�k�^kjl�ѣ��!yfq#��c���;0k�eBn���������0�Y�i�sc��	�~�O�S���q�`���/����	4 ���c)�A�:�,�K�i,��!'<7���K/��[�f�JJ�~>��y���&m���H>�b�>3�̒~�c����=v�1Ǹ<�e��+�ro�]^���������2�f�s�ړYG�R=}�Nm�|`F��2��A�o�{���� Y�A? �a  K�2f��3��t�-y��ѫ��=���J3>�~���������Vܳ��@Nv�`]�~]sYY�O��'�q���y���!C�>6l�П��8a¸��-	S23���z�O=q�޽{���e�vw�� ����|�42��:8 �����O���b�1H?L7��"�����@�~{ "#'Ƌη�p!`~��<ƃAI��APuT�F�����
� ���#���!³l?WBW�K<�<'x>J���:�&�S�W� .#�	�K���"�{p��q)�s��sP@����®�+V�L��j2IL����4c�6�P���V\f��p��H��*�eEC
m��#�b���K�f��l�KN���s��j�u6�Xnz���9:I2 � ���0}&i���2�Z��*�\�<��̜'���@�-C���fZJR��AaK󙿔�n)�2 d$ut�H��f�m6wB��etYvo���j��\�I~��J	V��?K8ȑ!�l���h)*_xNZz�msU�mm������-ն6v[}׀��H�+wȁ�<(�[�����t�b_XQY���> �
MF�vじ�������7h� � !`0,~�1�j�2�P_�1R�X ��KZ���[i;�H�(^IY�u�vXc3��m��2;��\�\,�t����駞�:�}����_��?Z���SGϠ
%�M�O��o�5x�ϡ]��
倥r̠��r,)c�|�����2L�X�ф������X�DYĳ��/	|K�h;�!˩S��b�e��YN��3���.��s��0B���P?d3g�c62�����7����2���U9X�P���<g�������4��B<ڞzC���:������Z@�i��-���ܜW;m��-*S����x�,�̌\��l��GH��$���Kp���o#���iSw	<q|�Rwp�o�J��g�Y�<���V�mo}(��F�R��̳�2xMd�[Yy�e���J�1�L@H!��4k�t���w��WH;97�m�U�~�A����Q����#ڂ�c�P�0���F:F%�����
����	u��`��t#s���q-D ����s�r��������{ʾe�f�qc/48�,+#A�9���AV���>�냻}�	KB�?w饋|����..�%��H'��iR����9f_Am�� ��D?���7���E��5�q��$�wB�vo� M�E�� �$�^�b�Xr��� � kd��T�{�|���ӥ.��������FbH��?3PFBb����sxf�����ϗn���[>r��ߜ1}ڋi��;�n��q{N:���yy���՞���TP��WTT���奖_�gE��~�7���ۓ�"H�g�Ո��(�m���:�u�M]]]�0% 31(�4: G"|+8@�
ܳ�h(q�$v��e e:q��0
6��N:����N��,9�+��M�%w��a� �Tپ�"]��{�S�ID�dI�#*�L�1���'
𠼄�fʋ�G�.���g9�=	�F�)�� ���\��/ e�?�_=�A�!b����4ݣ�aD�H�����HqJq�g���d���X�~)F
%��v���6qH����p_�����ZH��}0L�[y���6����v�a�a=�=2섶~Yj�}��2�C��B�g;��Z[�V����$�5Xw�^+����K�`���b����>u
=^��>)�Y6 C���u���L�/�i2ݺz����:2�Y�w�dYw�%fd��e�C� 8���+�}2�5;v�~���adPm=H�������gaMy�wO ��7�ͳ܍��"�6�����JKʬbH��S���yGډ'�h9y9��a����P�%6n�)x�ݕ2.�Q<q$Q���\�^6F(Q�:�h{����#�+�b��&#�TJ�+����'~��e�b��<xN���L���p�8�Kg�}P��qe
�B�`����p�h�w��i*�ȓ@̟���X��61,����W儯1
��F
���;H�g��=+��H!Ǜ$�R�H3���C��}ܺc(0�M���ŀA���= �AKQVB���z>���c 2��u"�zF�w�u�3�M��-M��X����OXh�'��Y���<;��]Ѭ�kR�v���>+4s��Ν;�&M�be%�>����3��d��JLm��	���"���.������A�����C�2CĲOp.(��J+�|ee�-_�����x�\NY�0r�����a��Վ�cF8�Cځ���"�#壝���Ns��>�I�9q@Ql�D���3�����}��">�F~9��3-�#�D���U�zt�*_�L�3���*6%�9J�+}����ghH���C�/�uEn�Lh���l���̦Ѿ^F�����@��:��Tr�A5p���e��!Cw��$>x�=h�/~���o}ˮ��z��+��������5.����� ͒_���`v��%=g�Qv�g�e�]�K���:}�6�R�BqQI}zZ����~��Sb=i�D �	���a�k�������\~�e�w�o�������_���u$�A������G�F���$IEL4V�2�۩�m��@vvf����۶mQ���V��<�wׇ��e
�ic��9P�Q�!��2:B@9"����p%!*�0=��ChE�'sB�#a��Qo��3������H�C����,"%�nkmk����ڎ][T�+*ͷܢlkjo��{����!%r��7V[��XU�[̣����UA�HKS٤�g���L�3qj���f�����p��i(�0��B(��-E$'��ڥ��T+���}�����Hi�.�"��20ok������:*IH鵎�f	�6�,��dӇ'ٰ�6+�PH�|}��!\�I��O��i�ؒj/on�=M���ds�ڬQC�]����r02����E)����w<�E�@cDj@G��k�
��Zoݭ*G��u�?in�X�:Z���Y92B1�Bƴ�7��,�&]��Tseg��@�u_��u6�i#
m�h�}�Kk�z��QgYI�����J.Ts���|�ִ��7�{)0�>��Wg�Yg)���a���)�%�2E4i��)��ON_j/�F�RD}�f�2)��v�E'I�I�h�N	�N��Ai�B�kT�`�b��N�+�gT:PPG�%ƸBi�}�A\�o߾սV+��s��1�h�����gؼ�C�9���욫��s�>G���=�N?�T������J9�L
�>��+,ȶk���~�������s�Yv����æ��I�������U˭���i I���#��B��2'��S�P�TOl^�(�2[]�e���;�!ݗU��xNJʰ��NR���5�H��Oj���Dr�R����0��,�8Exd� ��!��׭^o�?��M��Ν��mA���y��q���eJ�MxYj6��z�Y!�l�:�ͪ�nW�'���(5����@�!'8З�ő��۴��\Q�BΠ8�}!(�UU�nP�S��$�,{Ȩ��g?����𜶁��|�^ �c)�kO=��2І�,��ܔ�{�]����Ⱦ��N;�N;�t;���|X����;������킋γ�O;ю?�8�����#m���2d����Ϝn'�[�q���5=tӈ1��d�Ǎ���"[�~��ː�&e�����A^�����zz��"y#����G���Y��v�Z��'C��lӭr�.۾q��JI�jm��z۷c��޺Sr��2�3����6o��X:�������Nΰᣊ
-'7xT�U�Ƌmj����I��ό�%����D��0.�
VF0(6�|�egf��Ϧ�z��e �3�:��;�e�����R�Do�/{{w�����=�9?�2�u�qFI�0�hM��-���N�k�D��xJ��/�~�h���~)�-���t��߹s�56ԋ'P�%�3���Y�&Y�s�7x����J��k�'$�v�Wރ͏|���3R�M�za���Q�a�g�vIg�z�|�=e���Jē�Q�^�z�؃�e-͝�oo��/.*�o}�;n!����A�Ϻ����ěnz��r��6�p�O�ù;%7�q,�t}$3�������F����S���#gڂ������E�8��s�U�������k���V߰��=cƴ�ҧ��=T_�~l��w��!���-�����	����ѽ/��,w<Ã`*�N��*�:���^���ss�F���*�c��i��t��n$_�� �<��^8�DH���u�W�6�cAFH�������uLU#�d�a���WUJ)���d9$!̈	n^���kr)d��+#�qi��E�0]dD�#���(�sa���$���9Q��܈	���Կ��o�o�����G?��|�+v����fؽ{��u���:	�ru8\|���~־����7����'>.�t�A{��v������=g��eS�F�}��ϗ��<�E�cm����RV�m��L�={�ee���lu��c�
~����%f @�*�fn$N�8�f�n�'��QFۉǏ�#f��^+�n���)V*��d��P��\�:�vV�e3'����	�n�>�	�)3��P�r���^)�߁r�`��\R9�'�I�1�4ԈW~�~|�B�~,F�����j����>��&ͷ�"��Xs}���^�W�P��k�i�ܲ�
��ll~���fGO̵����1SG��b)�R
}�"�[�d���3{'���<�)x�R'�2:h��c���^�K4�}0lB2��D��n�i{�.\h�/]�~a���2���7�k_����я�'J���-W�✝�ae��v�UW���_ms�̴#�L�w��B���+��3����:�.��B�5�pu�Wk�w�[6oq%y޼�6w�R���ʻw��#<�mپ����a#�׿�u�壷؏�c�7:}ڇ:��;m�l�q�!;VC]��qp�Y�0+�'���IG~�lm��G:䉡1j�h�P��缧n��w��Rs�,\#-�'�o	|CH��9ˋ8;����UU���3`R�{%H��38da�����e��������V*t�aų����ee�{�ai�e�#x�?P���L���= �Q@��t��w��g���/�W^2�"���L����r�G�2�9��ay\��	��y�](Cn��I�15�.��";��s�G/8RF�7�&M� �8��/�k'�r��w����K.�K/{�-Zt��q�i2Ƨڐ�2�rWءD�qW�TKN��̘�.�!1P�Cá�ho|�$�`f��`�72�Ym�K���)\�a��\�?��sz�isf�r�����8���6m�h˖-S��6u�d�l�ĉ>�E�1p��ūF�J�3�̞F���HQ١��Æ���H�(��1�9�~g0�Y��:�-M��(3(�i0��Lc,{℅�#�8�1e|3\�⻰&Վ�7�g����"��`�����d���S,�}:e�.B��j�@l��O1#	nv���ZZ�;�u�?����C��Bu`I-����}��%��V]X�H��&^~~�m�A~���;���⅃�_x�y?��0���	w�, /��5��t҉v�Ygڅ^�.�?���5�y��]�����_���&������Y3gn>�6J��F�3HI�%!�"^c;'�6�HQ����ϸ�
��޵����t��_�t����q�o�f}�/��]��/��)X���:����tWWG�-U���b��%�+~2a�'q%)�sU�K��w��K7O�;$^*q�'��sLK�ؠ7!>���Q��q��<#�������+�t�X?�y��� yp�����c޺ߒ6���ʕ`n��鞱z���tuu_PP�F���<Wd~�ag`���;v6� z*�gAđI:F=Q��1�>�[e�|�AX<�����Qv�	�I��l�>��o0�ԧ>eǩ���ۺu�܅������믯���C��ww�I��ܳϳ~�v�Qs�P+�����v�O�s�����p�ukU�^;���������s<�뿾kw�u��(NI�Pu�u����e9EŶ���f�|��u�ɖ*C�w�wۊ5��+�df��R��K
zR��Lw��^��ʔR�6`�L�˰��i=�;f�H"â�'��a<�z[��u%�8�_Z]����2���đ�v�q3��r�u6n����� x��>���A�@��׫���[�ӟt7���e�Dhc����g��g��^����\8��JT�:���+�4�d�e�[_�{y�=�B�mm�r�e6t��4�_��hw��v�Yi�p;��2�Z.�Fi���m/���u]����X��^�DO8��@)) A�oڀ̤^$�_�{��w�6Zvg�]s�d�]�m7^u��]��F�P���}�lѥ��������j�O�H;4<\J4Mg-��<Bgy�{��痰�K�?a/�����i�XӊdJɈ��#�2u�P_��u?t����Ӓ�3mߞ*[�j�+�(�(،���.,)��;�h�S&�Ee��6�t���^?��G�=WfS!�H3ԙ�Sg~�Q�XXzH�č�s���bG��פ�"d�3f����kKm˶�xD#���}#�������tc�H�+�|TQ��9{�����+��=��i�3-,�ݼ���
�%v���eOu*�ڱC�I��5ە�ח���bIKo0������L�y4l���78c_�c�
=�[p��]A��_��tQ<Q�I�ˇO;�T�7�=�z꩒i���K�@��+�n��?z9�:�,�y���C60�UPXl�-��W�Q��P����<P;$;�z��O�xZ�}�ԟ��!��[� �A=�_�ۛ��;n�w^~��{��d�]*��M��k���K�q�t�9SF��;l�(G��VK�\n]x��s�s�6_Z<|��z��^��^9��.��ݱ}����{t�#j����N��ϻ����?�B{�����[��7� �tQ�U�����7�G���ʲ�#��`!Fn��d0QH�)}����[E��쩧���6��8��6o٤>�Ǿ����{��A�W��7���]-Y�'�Va�Y�2�y=�$�p(�J��-��\���X/��Ʀ;l��nd�g�����}ছ�N�g��MR&��]9�f��9�A�'�!��P,q��X���s�ۘ�c��sγ}{+�ӟ��=��S*c��*8�xc]��n!e��Ơ!4(9�ʑ#u������M?�~��ߺ�t����2��KnYz�3�F��%�6"�iC��V�tc2�ԓz���� �E��EO��Г`��~�I�h��ewj�͙3���ӧ?�|�}�e�;����O�8��W_������wڣz#���z�_��y��$�x�o�-���Y����WkgΚ��;��S�L9���o���V\��_�l�jҤI��0���WФz�0��w��e_���{��7�6��_�#F�s��(���[�Qʄ�L�tu.LE`�`X�tt��A��
(< ��^�u�$)M�U?����<�wi�NV�~!��w���j�Y����$ˣg����B��g�yw��[�r)���{=OW�|CZ(��חoD=J���'��,��R'D�eЦ`�Q>p�"�L#�;�u�ĉs����0�{(�q!�c�v���!tUgB�S
��~�q��s>H���!S�0��脭���0�̈́af*�֮]�'���w*ހ��w�����X��A1DB#�M$��[wڭ��=���n,]u���yܮ�^���o���̧%S]�
G�}�3����'�L�'�]���ާ��]�|�)�MR�z켳O�ܢ"��<;��ˬb�0kh�e�[���e پ��IjꎬGM*sH���E��B-���#�s�ֿ���^~Q�e�'Y��^����+,Wz��	e6vZ����>�٪+�����u�(;aB�5��jmU2��,-=�q�wm��ʗ�N��+۟��g��3�(��{w����2�Α��yW���h �Y���<�4�[
�j���b9CFXu_�=�L��V�d�f��)v�a#���l��dk���U�c�=���e��WڣO�f+��X��96L�l�R���^a�o�1!*/)��K�+�du�,�� ��Q���w�K��l�����ݨQ��?��j����7�w��m�V�~�y[�En���O���Sz�nE��^��8�P�'N;�?~�{~���k�p���D;w�_x�|�A���Z���b.��o|��<���'��_���7j��E�e.��iƶ*Z����;���G��ԅ������'����` ��� ����Y+~3���G�j14�H���P�wJ	ō<�ȟ�pO>�#yD	�e׼�f|(k�W���W�%�6YB�љ�f�2��m�v��\a�w�Yu5{�gþ�t)#��bf˶l�*Y�K�I>���,Ek��C^w�W�_�u�<�
@�
�L](���m풝�nl��@1����a��g�0���bf*�9�]���uW�YnT[���)YE�c|2��=*���[��d@T�p�/(���xݢ%f�#�>�M"$
�A�����_��}����r�L�=�FH�Hc�["Ķ�~H�ë1���v�;��8O>��]r���_�HI)��ս6f�H��T�Ku�~
mӦ�N;0�'����v۔��e�?�7t��Ëu�,�8�V�Xm�=�������ϲ����v�)gyܺ�F���K���R;r�L��~���+���[d�/Zt��X���s�I'������w:�ዑ��)�Ѯ,G�Y	~��B�s�n[�v����?.�K��u��ח*�N��W�l7}��*y���6��k�G��3	z��M�3�m���fY��𸣕�(�-EFP��9{׻���!�[�m�w]y���d���a�>EƜ�N��	���]Ҏퟘ��<��Ѐ�C	�ˑ÷��Q�O-�~ڙަ��>������M"�4!���4�B}�������������\�@��$�+:_J�tv��Le_)�L�'��'�L����-=�<�Rv��qO M�4��xPH�VD�*��d,�c�~�k�����\���������Mᙧ��}�5�����w>�~(/tGy�`;�Ĳ���м���X�H7�78g����]_|�����/�����@z���������\a��6EוN��+_���^{���@�@Hݱc�P	��R~�(�㪫��I)b2E8�*H�J}M2�>� B�$B�XI�q�=HT'Έ��a��Doi��� �[��[�N��%�3�!`0.eIRzIJ���=*p  ��IDAT�s�q7+���:)_\k{c�>�qϕ�b��p ���{� �.��y�7@���0JE�faa!8I��e0Z]YUm���YB�r�
��ÆH�E�Y��R�X��8���O��o/�t�9D�����ۑQ!�!�J$�P*֮]%�a���$p���/��#(��G� (�{��S��C+��*ӝ�����{�>��K�����w��gY����锂�j�}UUv�7�������xcx���J�]�~�]w��l��R\Za]ݖ��o�.:߆�ik�Z�t���)���ZK����$\�)�?Ϧ[V��z��m@�;e UF�:)1|�L'�϶�4�k��o}�ZJ^��J v��d��˱�l�Q�F��㭻'��on�uR3
��cG�ȴn�hj��Kf�>�M�e� Ҕ+a�y�p���������Sx%ep�ڳ�iÇ�/����8�4��7��J^t�Pe_���!��շ�K�U>M��S`�ic������ڭ��Bu��J�='���y=��ӛ��+�r�&�oi��*�T��yV:o��=�$���VFp\@�O8��@bɦ�a)�i��Շ�>�A$�vڐ�N;}z��x�~������+���͍2���G?�1�җ��uK/������EV_Wk�|I^�-� �>#N�k����3�=r�(�]<S�#�,5�S����k�7���t[��e��6m�$�iv����f��|�mް��q��)�����7����%焁�'�zt<A������̻����샲���oҁ����*����^g�0Ō!������5�DA# �
�KPr�'�W����},O�w��9Ʒ�,����	t��v�3�\&$i[���%S�ƌp���2c��=���)����S<��R�J}�Զm�}����B���%��>c��Q����0�K@(@������g�}����?��K�J%���,LO�1jQ�²?GxP��~�S���������}�����(c ���N�1�Ǭ7�)�G?��l����~���x��>�h7��O	0;��_��>����Xo�q�1���j�+Ғӑ ��&�K�C�����m����~Ϯz׍���ǟ�K/�ܚ[l�
�#��%�^�	�q /��X���`$�d�?���CXR����2L�;�����$�dٚ5�U�`ZFf���_ع�\�y����ˮ��O<jEH���_�����k����ۅ��տ.��Cʽ]0N�38A>��va�>�
�J�
0����hj���Z��go�%�U�eCܱ�3K�կ}��R�Az����{���o��L�%�b�2-��C\� :@ſ^M�,jhE�M�8�Xar�Y���9�l����,�m����I��w�#�Br*��@R0�V��*��| �@W�v�P^��T;�^w��VS����c�^��;���R�y�{wx��"I�`� �n ���ǰ���J�J�ӟ��M�0����}��O�V�*�b�C
9I�d�}hO��?r
9��tpJy�Rx�k����=���^�?Q���绛n��}�c������W\I^���?�n����oO.~��ko��{}�}��z�Ԉ���F|�� �ŕ|��iD�| 4��y�%�����vl߾���}��d4?;���˗./�@�̿RzR�Ox�*��nC��7K��/���W�z��W?����f� \p�C}���d�,e�<Ux���h	�R�����<���5[��UVV�)a�9f̘]3�,���(�%b�O��OU�Tݧ����J�H�@��<'�:�4U���<AD���R/E
y��&�Y��%+�_��U!I�&�:z=w� ���������k��ɤ�U��{�V�����E �C��Ԑ��{~�.�IF��;~ˈ2��M|�Ѡb�$�
=K�X��i�fkh���ԩ��//x?b�^�$ߤXoK0<�%N�08KKP2 �@L@$��q�w�)�>t޸Qe�٢{���7&<�2p������(�w�q�R8a��#B��J��쥗�������������z��g��Cp��,A�p�2���OYsc�:�l�����ά�_�����|�3R�^%�l�i6T�>u>YE��Wj�V��=��,#;�f�g����5u���cɩ��� =���nD0#�ʵ������HS���!������ӕb͝)VӬθ��R��(��ڜ�v��b��m���q%tU��� X������ꖕ���_����w\bZe���W�޸�?�<�A-������N ����ff��>S�g��K�Ȓ"<r�h˔�b{�5�g�V[��6,]��c�= �,��߳����M6��J �*HDĊ�
*b�ػ"���j�PCIH'����f{���9�Y"���{������S��9u��{u�b{ꁹ�u��k���.C?>�,U����-�(4�ڄs�eW�A��k�QƸ �XΑ��N��x��]���c�~�0^\d�<��+k�����z;r�L;��Au�;vy�q8S8�`0L�p��yF_��ث�L+{V._io���͝;�O��W��{��=����9~�L���R�3�}�}�-Y��}�q{��矓�~�϶!��32���^���� � ZĎ&'P��MVk�["���#1~!��n�D��>��G2��oﾄ��efF�'>�2і��}����QW���)7���L���P7�����M��8�;jG���=�'���De�7�|��75���荸���Pd��+���	���&1�f��<h��	�E8w�m��ϴ<��� �ɩ��n2f;LJ���1��|\�3��
3ND($8��G�.6K/���q�� ���/��s����M��W���B��0��;ݥ�W��;�^x��͛'\}�'�8�n�p����J�E,�5kV���"���?����׿�zǌ�}��8E�A
c���8F�1���!%�+s8�m�ĩ�|��]��'UW���%&�Y��vxU2��8͘q�������(Vt�l�,��Q
�AA}o�j{���WJ�f�۩��dcư��TG�h�!�1Τ����u�8D���󕿱cG�xp��@^�;���'�EN�޵SJ�.ۻg�mX��ed��%8S_��LB�0�$�o��~
��S�=��c�u�&��A��J&\�6�hcp���V.�&b�f��=;~��2�8 X4'#�/^��x���Q�X9�0�$)�ջ�@� ?��/��,���G�F���9�����d����ve��'*��}.�U��E�st�����̌l�|����z
|�zhc3J������:x?儉c��VգO���x�̠,�}	��9��	=�,c�=t��W\n�&O��k���=\|v����ȝw�1�I�~��ų�z�tH���:��|H
p�g�;4}�o�3�Hch���&< �i�|�o�N�u����]'�|�S�������/\�2{��Ļ�J������i%�5�b��;�N<���z���T�:�$�!S�LS�cd𔔖��h�c�$��I��3�A��9H� 
WMc|��û$ �r�n�G9!��ɁHjO�O
�ʥ��|�S��������^�FD(;��;\)������C9��:H�O��#($�9�QؘE�W��Pg&�<i�$gf�QYJ��-@�ayw,�<���C�Y��ү��x�w�)�/m&3�������ԓOH���#��ŋ�w����h��x��ʨ{������a�� �ү23�p=�f?��]}�U��ko��R�S\f�vns�3C3f��$��Ǐ36��_����/A�kg~�L(A�(A˘��u�op�i�qӧ�@4l�����)cm���K��v5ZLb�u�8N��::�����T׫�D3c���1Vz��1В���$�jh���Fk�'��:�\�)����Z~:�6;��<Q��J
�G���0'
�=(M|�e���%3���3��>�1c���1c�q6n�D�I��d),�l��1�m��i6a�$++̶�Cr�$[��Xm��_���ek7ڂ������ *���B��.0�ͷ��\K-+���\������I����#Y�[���|0���&R��}�~򫻤��_��Q���)$�D�PB�
�I�n���3Ɠ��|r��eRj���U�`�rs�`�O�����4:c��\���l��ᖗ[(<��\_�ݹc����}��E�,J��~�;��;N�ԋ��ڊA�YM�8�N����R���im�h���;���̳C3؁�?B�o��u�W��O�"G��� �	�s��E�
�p���h\#>H
<�w�Ȥ�)�E
e��5����*ľpC���J�a�>�'x�8o�JH�FW�pMe���l2�F&�V�����<$�Za��E���^ڃE�_�Lho�$h0R�#���1�y�7��aq%T{��Ë� e˗/��.�ئO��#���ؙv�9����_���>>�=<x��ER�����΃�D���<��W����z^v�|%�+_�¾��o��ȜQ�;������F��:�5��	���QRR(�o	�M]�� ��/��r����U�^k|��������E��+W����C���ﰯ]s�]���G�/��}��W{��˾x��)�E��&�$�r�J	z��2a�-�����c�ɐ��!�q�B��LXB/�ȟ;�%߻���Dʜ矷g�y�'V��K�,v���cV�XY��K���n����&�n�?J�>~zZ�����@N��9�@�&G��T��!nD�d(�g�nQw�� G�w٪�"�Q�Td�w޹~@�-���+���:������(uPN����W82)��>F|+*�{�~<��ݠs��O�}�Ph�
Y�*!�V��B�=����M=d��V &<���~�-|w��#�*�]����í��$8ⱄw��i���f���)�n�E��/�� �N�9�UQ��C0��7��/��PO�D{H=mrO�Ў�L�P.'�#dH֠&�  �s_0��
�g0�]'+�J�}f!V�'�߼�e�o���t���;�Q.Wޥ>����a�3�+<�<����wy�w����KX��k�?��t���6��o *�Ih7D�[�WV`����z6��=��������=z�_�Pv{���+W��ݖ-�V{0c�A���^���C�%��Dݫ���|mn�qMT���AiE� ��%�H5�g��-�ƴ��m���V�~���V��9Q]��9%E��hR�P�'���NRg\qc�kH����I��v���u�<J�M�<�g��c�7,F��_�S�cCF���H����U�3�.��5~fQ�<���~�S70a?8����b㎘fS��i�N8���:`�x+1�2�s�Se�'�YGw��&٤Q�L�l�P�w��h��{�L��'�o,�'L�I�'��s?u�1��h�ƙ3nR0q�<�q�hi���B�V�د�̕�rUe�����~�F{���9���gۃ�̶���Ov�7o�[��M+߸ҊRS�S��P(`�C�Y���,C0N�[b���@�c��ngaCƍ��N�R�}�OcɌ
�f��q���A7��������<����ȟ��x���	N�G>		����6�Ey�]R����"���6�(�+���qhq��B�ϫ��TFSKO��բ�:�iEt�,��R#�Ӳs3� ?�W�r�	u��k�e�;V�?�⨭��Fo�-t��6��}Rho�M�/;%���2�F��}V�He�=̐�ܹ�yJe���>fyq�e����K�u��	�#l�A�����	mz��=�w�^�0"���n8����qè�5�U�f���k&jdE)D9�<�K9L�@;6n��x����YOU�6h��	��C�N�c\�x=��O{�_{��xN�װb�?U��U��c�L��p���E3�5�c�ʜw�*�^�1�`�-�U�A�ۄ�]y���<D�q�d��UU�?"�b�&s�<Fn��B�3��p�qa|�x��1.<C&��'��}����)(�ܥl�F0��J��#,E���wߵW�<os�<g���k��ܾ�6o�n�/U{5��֠q�����,�>}��ᲄU�R%?B��q)�f����;��ȿ 7Q�q{d�w].���$���#d��p%�K�b\t�'�l�OBP.�q�!���W����?J��H��Y��i�2�^����o�h�B���2��G�|���A�?��z1��c��0q����"�E���O�-�2Əog�q���k�w� /�������ķNW�\�$���;�M���Y��H�8��ܥ���[p]����`R�	id2�����h�P�&/�r�
�ͽ\�D���w�]x�v��wx�$������O��ֶ�ض���h�?���3� k�)�'<'G�=��2�<fLzƟ=���NR�*���F��&�~�-N\��������
m����1�F�hL�M�0��p�8���^oB�J��@%HB�l�|�{\!R@��@ܤ����'*;2 ȼڂ�����I�<�Od��.��ɤP�@l����.bŸ�oޥM(���7���&�������!N�#�D�A�A�ٽk�+3(o��D��O���$���҆C�'��}�.��EF��sgHFQ�3CD���͊���/��#1"b��W���i�9��vlۡ>�=���=��UR��E�6V�HK�,��}6r�S�0�d�0M;������ݿ�Z��iiy�z�n���r��ע���Dw��P��	�n���Y!\�0��+e��V�:c�,�$�Lf�O8܎>�X7}��d�Z��/�>�9�F,�����/��~Ŗ�!�K�q�,��l<PTq!Y�n��_��~�a��}q�����b�ņ� �"uݵ_s�|��h�~����/�M����;����ϱ��9WB[�?u�}���ڗ��}w��)F�П���}V���0k���.�e�XV��6x��x��6��Y6x�8˔�ۙ�`MbF5RH�w���N��a���$u�#:�\quc�@	%K�������K���2J(���>��$��}�0�9u9n�>�>BP����V]U㊳�=��"�r�j[��=��(�:��-��0���%t0W�6SOx��ׯ��"�J�)Β���$���$e���g�@@w��7���W���2�>�rx2>��9W��x�o�} ���C��d���&���>خ���;��g!�o�<'���{��^��}��邺Y!�������;#����f�3�=�P'���JVS���[6���qe�U�$���}'&L��(�[cG�^�&�+�� W`���1��o{6w�-�ʁ����q�G��#KhJ9<��.�-�E(봉q"3�F໔%�pܦ|2��.�� �x��&���M�O��'���GK�b�46jC�_햟�c#dP��dےŋ췿����|U�W^���9s^���x���g��\s�{��}�Y{��g�{�g�n�p!j7g0E�5Y�YQ�J��������C�Y�c��+��ڝr�6y�4;�����OvCz�)v�����2�?v���z���Yg�m�s�+�(ߌ#�����p$}�pX��+���A\�g	��И`1aF�뒒>n�ڞ�:h �\�֮Y���}{9-2`�8�XS&��JoƝ>a`��``�lJԷ�<��}u����m?T��G�q��� ���K=�����顇��Y
4����ϰ7�ě��0\h#��ƀ�q08$��=�X�<2l��fƍI�#��c�+�{LR�<�,�Sl�c�����%��I��x��3.>>R|�A:PQ���Ԙ	��/�p�+1�q�P<d������~'�m���7r��M�����%���W�ፚ9��g҇B^��I �RUU�lպu*�,YV�|���;v5�ر�m۶�Tv�����$���� ��ށ`bդ���9�w����߱Q��[~��<�g�]�����g����f֐+e�\W�ja auގ�V����0��C�dVr�Ji�O�=Ĺ	���V�`z�Ƙ�`�(�����"c�pE)A(�{�W�ڢ�u��M�E�޽�]�kI��/b�b%�X� ga�[\����;�;0���jaN4띐Ȓz�r�&3�Ѿ�� p�u���gE	�k\��Ā`�X�>]��&1�5b��*��ۺۥ����Y��65���?}�]s�w,;/�֮].�nQ{�lذ�bT�ኤ�j_Q9��sY�՗W_{�Z�WV�h#�Gdyꗛa�-�l	?�K��R����� ����;��ږ��om��2e�j�%tH�vJ�Կn�)��dcPh�[:�LS�i�V)\��^V*8t�F_�YN��4	��FKM�P�^�k�v�}�����z�]����/\k����K>k���%v���g�gg�qN��<�>���_l����r�:�1�H�W������{v�,3{3RR��,����^z�U	�'u}EB�]{{���p�2[�r����c�.��7��qJKOsϷ�>e�]Pf��֕�h������,?!�:�e��S
,'�����ﯩ��&)ԝ�V��j݉RN�3R�[%��ڥ������(���461R���A99э����˭+)�bS����[7��}��܍C���oH�à�q��ǃL�b�?����dy�
$(�	���+���4K��S�b-%>�bUn��JGєB��.A҅��7���
�z��X�l3����$�#Z���#C�	)©�dxR@�#��Y0v��y��w�o9���ߑ���B�W�Y�'󻣝�7&��� �*Y��ėi_Ge'�}RXb�EMv�#4��m�"㊒J����I\�=�ⓥ�X�ƛ��0n�WZ˻�~K�����I�ňn	� <��dA�=���B�x&T4p,.)�i�'���}-6��Z�묽�����2�TA6X�g�х�چ�<���^z�]�p��9����⯜�/��-��M}ip�K���M��(r"
 ���J�0�C����]Y]�h���kØ�U�pY����(`��E��/)������A�[�t�-_��6��l[�lw���w���n+ޓ��t��^��e3��+4Bۃ��ϑ9\Q���MVؐA�;��?��+�!a �~�%�7)���*�����:;d�+��83V���KK��S���4�FmG̜e#��8� ;?�F�k��u�]29N<,9-��o�$��MQ��E��m� �G���C��Q ��u �Cr����ډ[TT %��vl�,�8�&M��{dje���H ��^�[N`�;PYk�6��k6؊k��n׮�p�d�� �)����U�5x�K�͊5m�d�;��dH��� Op+㻢"ܱ�WV�Z,-%���l�v�K��7��S�e��ظQ�-?G�<3Ǌ
�������!���\1��1or��"#3ՒS0D�Mx{SeH��X��0�;vl�l�Q[�m��5�]k}J�d`ewRe�E8	�)����	Z
�N�((�u�����%�B��~������{�e&�Ǭ8��[�gL8��������Ŷp�R[�h�-ҕ���n��w�~����KT�B'��wY�$���: �,^'kd�]o��͙5�5Q8��֮_Y��֒�|�	�y;�I��������q���M�^x���D�6� �9M)�.��흝i[�m+���9��1�w��
�ꊡ��me�9ף�
�c��?��H	�<)��RP��X��u�����ٷo�61�)�YjX�]x%}&8H,�p��u4Z�ڄ��hpdR�w���7���ѵCV|���&!9a�SŸ�ET@�3��/��ԥ:�a���:�B?W�wT��<�ʘ2g)�o���=�����%$�����"2_LggG�����~R��[���i¥K�<ܷ~��#��V�7�n)$�2P�v�Ѭ{M�j�)r}e�Ŷ�7��R���0�p�S��sE��KB4�VA`mdfIX�gd�g\h0 |�M
c�A�wl�>���:�>�|&b�1c�2�WBpWd�4���R���.��.���g�!���슛��K?q�]v�E���7챇�~�^A�3�Y���wٷ�{����������}��[Y���}���w�,���?��J���o�m?�����K/���v饟���/.Xg[kc-q��RJ,)5�b�c��3Ϊ�����⥨�$�Y�r4��jW�m&]��Ct��x	�6)�-lD�K�fK�L|���#��dS��mZ`o��f����U($�}7���o�I"P8p���,J=Jߑ���݀���q�nz'�B�x\	ߣh�:�!��,#rGM���z����r�T�8���|�\�\�b�L�T	h��j�R�D����R
� f��e��Du�
�T�j[�ƤC0��0һbi�Z��#eaXa�ծ�g�<�{K騵l	b�oM����o_r�ot������]��3���^\�$�X������aw��?z��,��+f�:�fΜ)g�mܰQ���3�/�y�.Z�AR2%�2�(z����Bۆ�@�@75;IF2�$�e"�2V�"C<^c��!��w3��f����K+����<�~��N�*��_�;ma��kx?F�)��>1�چ@�/>6�'� ,�V�P�X�`��]��.�,���P/bB����TYȾb�2����~�yvhb��z�c��O��	o�M�}���A|���������;����">�$J4�I�[2�t�2���'���a�qg�GʤM�� b@Yc�W�t_���gU��~�۷�u�]g���o횫��O_z���裏z9(��FUWU�^O���K����\�_����g��7�C�f��O��֭^�I���>	�GY���ߖ.�
�G�=� � ��OƉ�|�}���W�1�q�ĸ�-���R���w��K�0�/<��]�ɋ�I�р}�UZjG0�V0`�}�ҫD�V_� V'�H4��i�dFA��=�
�fpC&�;�.�˾v��X�������l�����Ui��u�-��A�~������+��mۺ��;�[�x��7��oޟ?��O�-�g���.��9`�Q�1&L�_�)�?�n��-��[ ����޿:�a��߶�~��	��U�'.��]���yu�NwvaP"8�%�=�������8�n���-c΀'L�"/�X2���߈�B$w0"ط/]��$l�����@𼹙s�8r�$$9�&���'����6���������L6����8����?���S	��U�c2�G?��������.��2�E��/.�1���yh���~�w�_tL&�Ё���*�M�RԶ(xL�p�}Z!?|[0��dx4+R��ĵ�����}�9����V_א|�5�|��?�w爑�Si+��ӆް����Dy���J٠�Z�#>{�{��"=k��e�#G���C>x�t���U�߸1M�NPVv�t�� ��ƛ��}�ۄO��H.��v�w&iX�+/��)ZX$:���3�\���GJ	:�"� Qݺ�;^� Y��~���>IJxm���QBn���
�z���}2��3�v"MHh/..��v��U&D�>�K�*��a��Q���eR���r%�Y!�1^0�:�m�r��F���n7�x��8��9<�[2�Qz�Y�L��O�1�������z�'q���w ��W�|�!J��nW�����Pv)�ѥA�?\=8�%��'
ª�U�CL�
a�� f �Y�Ng�0��y�6���6�`(0�c	����;�N�{�GI���]��ƏW�?��$��jU�Ǝej0	c�λk�=���t���>f8j�J���F�@���.��>�	���x�!;|�t��?��v�W�R�[}���o˾�k�Mp��_����=�k��/<׎:�$��p��hH�����,%�%Xq�>�ޕl��*=��b�g�����2(����̶����O����D)E��&�/a"�@㓙!�A�� A���aG�b5K��k?�β��Z^�kN�$����B)��Yx�>c!E�$b�����2F����T
���}e%����H-RxC�\��}Q~j�=���]5�>�(+>��5h��z�8[�i����;�S6Rc��q�U�s�^mdEI#�/�Zt/Ie&i)3V��Փ;E"���<h�$5ƚ��wI�/J��=��~m-��X~N���d;P����}�����^J���ģ���~�gf�i` ���?rH<�����v����5��ګ�َ�;l@�VRRl��(�ј����]D��� ���g(��5z�I� ��VT�G�m���g�i����2a~�+�c�JOjJ��i�+Ռ�x�a���`\���[D��(n�����E�buw&����V_5�=c��w�9׷��M/3����j	8$�E���܋f��?�Fy׀��@:GI`�Jv� ��%E�r�w�#C�:���=./���EQvQ�}|G��I���hkm�r�!	�>
�Y-(*.�!���#����
��j��%�̜r���LJ0�8�u��_���u���s�7x &:��N��B�����٫B��H�~Sp�q����(�D�G�}�+ ���+�سk��3� �i���qm�_���?�D����'�	8R'��<'������}��;~C�R�9��{�O^t����s�_,|�u)��MU�7;�&N�R��c'�y������"�u�zL�����0�aιVLDp����j���mܼ�~s�S��;e4c =m#FM�1��;�s흅o�|5j�˲�'{�w�.���3O���R���9���6|�\�#J'	����p��'�ѣG؜9�iL��ꫮ���g7zX}���[��k���o{�V�@��O0b��Ǫ���$,��	n ��������[��'|E�F΃��>�u�/9Z5c�ȼ��A���.p�-�g<ø� �L��7�G4?�Vcy�=�ĸ�Vx/-5��brl:��Ν��]p&�&���z$� �"����;t��)}��V�X�Yd!U�Rn5�5�w8P}�&�S��h�`�Ì#2�g��*����$ʈ`�\;��e|`���K�Iѫx��/�<����!���6��+�r�����c�NTS�c�gR)���	��樂�{D���.
 �ÄD�����1hwl��"�Xp���t������#�=V|�]w�y�G����_{Yc	�� ����E_��(]XRR�2u���W�@zn�h���}�c+�㏘�g����?�D�"��;w�ZD}���}�|&��-��{�Q��Z���ۤ�0�D�`��,\1�`_�gр����	c@U�\'`H�����/������}F�p��َ>��1��%l?,�I�x��۾g������6iȨ���6m��FМ9���ߺپ##�gjEd�}�z���~�yḃ1�������ek�]m���v饟�cN:͞z}�m������uZy��?��ҳ�Zm����jI�)2�ҭ��U������:=�r��b��F�o�L��"�A&�S�Z-7SvmR��]��Rۚm֔���gm��o�������f�b�(�8Zts�Rs�y��'���=�
��
	�a��7���V�w(�ox��$Ǝ�=W��.����+Y���[��M�I�|ٶ7vZai�M�>�{i�ufZbF���4Z��8�#�?I�;�8�Q{\�5KYI�YA��U+E\�8Pwdd�0K���h�hi�Q�ٖU��^��V�m��e�Yfv�H�tW^u��s����G��\z��+�#Da$!p�5~A�� !��~�1AIly�J����AGye��t��O�~e�}��c�<᡼�W���u��^�Ɣp��APN�>C��ڛo�%!�1ӸS��ϭ��Y����ڣ�0Q��#}`�h?�DPf�k�&2�� �{g�HB�#�o�Š*.��-�����;}|e�Xf�G��F(�w�5�"P?�<�̐�|ݔ��	)�!c+>��|�5�`��v��� .2a�'S�7�W�=�2
��sf�7n��u��qGY!�+��
$�����ǉ�U7��w����\��|�
$�0`����/]n���������n��z;���-��g�E�����q�}��-
�=�������~�R=v����-�����.��Ѷ���i�R�	-��}��~._��v��k�}��G�[o���Cfx��7`G��;SG�<���l��{�����\�~�I�t(�sϼd������JJ-'?˒�1%iv��gZ}s�ն���,9f�7��s�ڭZ���W&D:�,)[�͊��?k���Zn�`�����+o.�������Gb<N���p�=��_�-g�}�1��'��w��y�^�ܜ7���=��4V����u2�L<�Ó���R2	x3.�)�q8���W^l��k_����㟝�SS��'?�ݾ�E�AR�5v�E��yo��}1��75�Ÿ��x�y��$����*Y�,��N����#0����h��oƏ�w5p֪�_�S�(��/1�
��'`�qڤnh��L�V$ε�7X)�𯷁���{4�Hԃ��?�鏭��X�罶a�&���3	�c�6�P���)� ���.��+���=p��Ʊ��w� ^8�2��c�u��>���I�����?��g��y�xH���N���/��_�zǄ�S�1f����x�D��X�O����l�Ȉd�"��l�0�@�/�]����㏿K���z�x�W��ּy}⢋�������¢���4���EW^y��*���aLi���פt�������g�y�{=������_&]u�U�?��O��;Ny���gϞ�<���.̖,Yj�.2���"�ɶl�b۶��ed6�zI 0fk�R���!�侙Rh!C'A���Qtxƙ �>9�5����/p�QGe�B����g�p��o�G�ۺ�Z?�~)?��Om��m~�Q�*XRj�=�;�Ɂ��R
֭�`������U{R=8C��S�͓�yϟ�Q�El9z�����C����}�v{n�)��6y�2b���Vn�2j��9̦Ϙd��ZAQ�ꋵ�V�G��X/!#�$^
��O[�%�Pb5	�N �fz�H�"N
3�Iq"��+�H���e������W
��m�{�ۖ���S[���N��	���H"#|�E`�$����C�1B��[��5|G9>v�H����s�DY��סk����ޤ��'Y}w�-Y���[�,13�dE�(��p���j������#Nj�1ݨ�Q��u�a�t���b�<c�Ջ���ݹ�6.~K�W���0Ϟ�&	���5��9�SYk�mp<�Oť��W�U f�,�|5����i�l�СnP�o�ns�1�\�4��8���ΘN[�n�-[�Z�)*��q�P��xK��M7��?~V�^�{P��YmU�5�(�δ6��8j�S�ћƗ�I0��A*||z����a��[�EO�]�&��+tL�1l�P2d���8WF3ٯ�R�B�s����;�� ���H@���` �v�ۣ���hv�o{�)���Q�����J����s��d��	<� f�9 �+��G�;#ާ�����O�{8t4��/��s��Y�����(����!���Q�0�"�Q��(O������x���_�֯]�]����M��'3��)9�ed�|đD�e�w�u�Q~f��ɓ|?�駟�
>x7i�D;���ċ���ӧ�8c��4v�)��,/7���&r�'��<��1��aLB��`9?\��ߑy�7�H��VjQ�9����8��:{����Kw���Xo�sR��#�8KtB���m����r�&۾�][��s�I�t׺Ŷ�wl���V�c��_��m]��M7�r��ymۮJPiv�ş��
c�I�r��m���NCɧ�z��U���Ȱ۫>�7�.��BWPz�a�[�/�>A""�<+x�&�5�Z���O����-_�n��b��q��6a|�z%���^��.{YR�;9|X��"8<����G�L�K�dL��>�v�>�h+L0v$�!×0@� M�x	]s?�ʒXbe�3��ʥ�6G ���ꚭ��E�#���g��^m�\�q����}�nEm�M�������j��~�aK�,s� Z�L��-��|�:i3�I
��J�Y�Eo)�1�6p�yD�wrTD�����«���*�=眧��O7��J7����_ziҊ�k�)�S�ޕ�y�%X����HVv�1�+s+�5ܣ��o��|t҄���K�-//��jԽ���ؖ�N:i�ɓ7�v�mQx�� }��O�ϙ3�x�c�!PSܑC{����*��Gy��?��� �;�K$8h��Q"�D����E}J|���O�I*�bd����¬!�&0Gd!�(AZ��Pa�(�G��&$�Al���FJE�+��e��G����� {�]��?�w�E�.��	<p�yv���ٷo�����k�y�0��?��]��_����o�l�����o��_a�|�{��G-5=��H~��_����\�u��_�C�r=n��W�}�;߶��u�}I�7�L�fo
~�mRZ���D0Ͷ_�w���6rd��ۻC:�}�x�[�L�~.�-9��Hq0��ٞ�
��'c�VE�y�͖k5��Vm}d(Ό��X�e �r4FJ7�b�$6��3&0?�5P�H`���F�`ȁ��Q���;�MY�3F2L��bk�u��(I�g2���D��`C"�\��M\B��8KJ��⬶�ъ
�,Y2�����Z�[�[Nt(�꟔��n���U��j�����Nu��  ���O�A7U����j)�2"�7>���y13�!�D�	���J\���U���=��}�+��,�{�K������U��HaY)<�g��{����#��;��Rb
dhͰ�O>I���=E8�W�n���[�nٶMJ���ĩS��/|�.�A9>�9�{���A)^�?��=����2���~�a��[�m���(��q';��$���#�w0��-V˘Y�wXB��_�4�H���;,٤^�P���:�YP���������(�3�2B�������hw(�ĸA(9���c�����0�h#�q]	Fq�.��F�	�L�	�Yx$�7���B�o��~;m!��~G��VeY=�q�}��;�ɸ�,��I���<���_������v���m����Oo/�Y����a��v���yv�e_��}��SG����=��拇�gP�Q@q�{�ŗ앹���?`���/�Ow��9{MC{	#�v�:�������3�����/a\��10��z��AIGQB1$0���փ�D�
	#�@��wZ����қ�k��6nh��(˶��f���a�M��/���f���wY�tV���n�*��aS���3X��Ӫ+�� A@��D���u=a�c��-V ���|���!mݲU���i'gh�|�B���� k���*���Gߧt�]w�~0��}.��m�[�%8RbR��Q����S۶��߾�7����M��|�^��s�>2�����|D��-�C�iC����M�+;���m��r����F�803�*�"��Du	V}�!Vđ}Y�9�����`�{����GH�MD�I��20�G�O�N����~u�w��+}�^H�<#9\����7�%t � 8���P�2&Љ�-ܧ=���U�l�h��"���A�x�?��>������y�]x'��� s~�?�%�������˧._�������$�����|�����I�v�c)7�)�zď��uk�ş���O�����N�kIL�C̈�Jq�����PgJx�dxru/ګ bB@ K�ӈB�"p����7�2�B�gYwޥʂ��]��=�`8���凨r�-��}��]��V,_a+���P�*C'��w�-�'e����m�����o?���{����y���{�+�s�YP�r������ʊ*?�_��W8���<Q��~�M۸y�+�6e&�YJZRJ��R����wZU%��:�t�A�R�ܳ'؀��2�DP.�\���mIq�i���FK�qT��n���lTI��+N�	ũ6sd�7)˦�H�,�C��ZKs���f��⬦��é��A��C�B�@�#J">�!�fø1~(��f��$ƌ�b|��}��i��(4<���k�}O�����	S�Æ��]?��*��2�;�8;y����	��D�'5��α������� )0�ݭ�!e$���Z�%D�,!Y�� �^
O[s��zI�puIXuI�p��q��*'�a���Qʳ`�~��l8JA��� ��}��~�� /��M�|Jx!�0232���.�YlJ��s�Hj����]�^�`�l�6��n�48\G��4��}v�]w�����8��6�T^~���)6i�8`��n��1܎�5��:�L;��m��G9]A߁����J�ݬz���ؐ�����R(1�=0 �Pd��Ø�l�����_���c�v)ĕ��.��q%S��Q��h�����_$����*^�F|q=��B��ʤM�K[C9a�h7�C�E#���Nx/�<(��hu�$���������{�:f����e�KC
B������`�1
}�y*������[�k�^{���?������O־z�W�K�	o�я~d����	������"mذ�/Yb�<7�n��v/�7�نM�����������׿�Q�+���'�|��@{�1���?�������k�y�����
h�2��7�x�� X�E�N�T�Z)��m2��{�X�p�b��������|���R}u#$d�Ƙ1�������/i�l�������2$�-7+�
sRm@i���kyY)�'?�J���s��8�2�{��륍1�)���]�E�q�7�@'��Uѐ���/Q2�k�o��c#���H�Lb``ql�'?�I��yDD���L�R��W5!�Q�#�F����8dW��.8���ڵ_s���}�������N>��9�\���L&r�/�\��!��A2�}��1ތ	�yI*B|�^|!�&M�d�s�q��Yg��+���0>1��F+�>��JKK�z9�,�sM>������I��G��H����M���{�G��W3�?�Y���^H>��cEuD�<��}2�-�Q��,�ox�ü���\�.\&�ä�٧��A������1���0
��s9cu���Ǐ}��[R^^^�u۶�W_}5��W_�f���$wk�F,�����	��!I�Э1���> ��k����,�@��!R<D��34�VbQ
�D8����O��2���%�!� 	�?~f̈���h( �����!d�/�Mo�&��,+nt��Y2frI0�.VmFI�spᰡ#m��Q�o��/,�Ո�jB�v�H*���F�ᒭ2Y��P�S��o7F���k}������Y�0[�A��H�Z)�%%��2':�3{IY�Mbh2RS2l�kmՊ�6l�p	�X[�r�o�OL�7,�C�tJ����6K�i�>٩6~X�1����e�86�N��kG��#���'X]E��UV[g+KX�>�e��7���%�p�2F�^7.}e�+
0G���LcI?|���Ŏ�7(<�W|�
)e����w�i������ﶻ%������{�W(R?��+V��կ�i?��v�׮��cGZeu��?�����5�Y��j�錵%9v���v��2;jB;jj_7���r� ��c�D�C�j#�}Ƭ��J;�
�g���`�;�G£3z�o�G�=���	Ŗ�&p��	.g�����w�Fh#8�/J
izF����n����W���K
QU��\KK�ܥ`w%���fXqS[�n�p(ɕ���l}��8[����^������<w�%�
J�~���[m������`k֭q�p?{���%1�A�c"�>�g��O7�7�EY��p����!Z�(���E
i^��������C]��h�ر�:2v�80e�d�{谡����c��c��rEĵ�w(��ߔO��D����*�E"�J�A9<WϽ<��;��
��S?u�J/Ϙ<�\����Sϻ����Q���f�#�>
Ly-R^R�xpQ����8�t�S�\p�z��7�oi�����U�����km��'�|�Q��{��6���g��|�~���w���馛��n�����no��/�%�6���D�o�<v����;��/�F��>�9�%��}����_���o:�w��a#4���;_��W�ʫ��+���N=�t�Y�p�	��Ҟ� {��t�P��'}�^r�|�֬��$��D[��-� �V���~�bL�R��v����AT��}��6�ԁJ�_H�;V���!�a�|u���l��� ��w��y��߄>�n�1���Y��3a��B�?�#��$ 9~�O�i)��׿�վ���ۧ/��}�������}�[�Ҙ�j�vj��쳟��].C;Ku3��)��ϑ�:� �{H�0c������}쁚<y�h �6o�`K�.�k��G�F3�c���9j�ԩ������8pN(�e�2��RW��n��� �/$�C���w~蜺����aby�^>\��|�cx��\��	��w(�J�vp����Eٔ��^(���uI�$,��?$	6q��5�*&���&��&��2���l�׹������w�u�)�_~����v�u�=�إ�ǥ=E��$�"�tj��1� �x^M]� x/�׫�H�_H"�X.ˇ�d�����Ʉ�y��\q$A��Brǹ"��ʷ����2@��><�B�<#�Pp3`֞�W�A3�m-�R�8�AF�T附W���`  1�ph��K��C�����Wڇb������>�H��-����x)-(�,����mRn�U��N?}���Ξ����=<&+�QJ*Q��D!I����R	v	�}�m�[��9m�3/��}������?f;7�����t%��3ϲ��s��:�h?+����]s�5��o�`���C���m������xϟ�?�����0���p��r)2a<��`���b�,�-߽Ů��������q���#f����]��x��i��V"�,77ǲ��-]J�����`-��-xn�B����'�y�^|��^�ݺ�-��Ί��mh%)W�����0�i� 7��o�w5)a��W�^8Fr��k�X��(���������4�
���|���	4�;��ωX���ۯ��J!NMϰ�������'�)����6J�e�
�L��)�'%$�g�++��y�Ǉ	g�Rq�cCQ�"7���(ޱk�+���5v>k-ڡ=D����BC��Їނ�> fn��L߹ڏ���B�s3�08��oi_7�(M(��B� ��HqbJqq���h�����|�j�$�vs&�!W�c2�����2�4Fa5����1r�&��6�F V�h
'eSWIi�"��{��c��� ?(>�Q��N%��������PLMK�ϔ�x���K�H�\�Ӏk��Ju�"^�Il�s��;�~N\	���/x�0*QX��}�ݐ�[�d����H�s�,R����QAa��;g2c�x���N��:t�e
���>�E���2�c���(:\�l�O�����o~þ����7^���9�x��?�o���d?��O��?���w�_�?����(�@����rIUՕ�/Qd=�qcOg������`��"��d`dhtt4[L�d���F��(6?*�$%ؾ�}�G�1z��4��Ao#�Ю�`�Y)�����O�T�yr9$\����b2 �:x+0�E�X��u�]T�5�#��h��+6Ӧ�c^�+$0�Q�g�)�ǎ�N8ޣ#w�qNC��H�.���v�W�ܲ����h�^η�З�Bϊ
<��A�-�/ܷ�������Bm<h�������+��+/�b����ހ��� � �=�˖-w܁Ψ�v� =t�CG���1�
�A�C�O���`~��7��?��aC�aU����̸D�Mt�r�}&|�g�p��6�;W��zTY�2�W��w�-ɰ.��v^uĪ|�b�u�=���5��?��*���W�������}��M��ض��?���|��}v���k��X]!��K+W��o���ɍ���hbtn[���e^n^�xy������#������t�7oJ|��7�����c���%�R\�@lz@8R�\�I��N h��~�zԀP�;vF�6����-6�NF���,!��

\^~��t�v�����!������*#֙gg�����%^��u��<A(01"�&�}�} <Jqk�A��ĕoH�o��)%f��[�Z�R�M�6�2

mGE�5��(������fu���-!)S�8���7�$��84^�p ��������^e[�o�/�as�{S�-[��r۸l�-zc��Y��j�ǄkK��z˰���#�og�q��r�Yv��2Xf��`�MQǏg�m�:HJ�`�߯XJl��II�/�6%9ў�=�WP�$f�xD ����!�eS�N�SN=�v��f�֯�M�D�޻_Bc�U�UZ{���T	��@)�R��+km��r[����W�ZuS���@���Y'Ť���w�M��ښm��~�n۸h���Pi��2�L�U8fz�q�HWb�O/WW��q�*\bb8p������d
�oX�����ι_���
�I'�$������c��B�*	<� �M� q�;3����;.�I\��D)bM�)��9��"��m�����'�"Mmh���:g��.�Vi���?�h;f�,�?p���X۴q��9�_Vj�m[K���ZR-M��n�d���4�K��@�|��/zp
fء	+4��Uw3�D�C Gd������a�z4���t2��@qƐ���=6T�3҉���b�^3��	$� ������*�i��ͺ�U[e��gU�\0gը�#��il��� ���Z����E������S��Єq�����<��>��TQ�*]�w�GD�A ��I({$x
���d�a��?�{��Lτ>a�9���c(4ܕ!&�PR��1�v\&��$xj���d9�i��-ř�&�����{2��k�]�c�0�Θ2T}du=�ƍ/�� �l�O<����{j�#���!�#�Oa_�+|!¢�Qբｻ�i����}�.pd�hj�ȅ��Xn_�`6�}Jo���ƾ�&N�h���l�f+V��k���>c����*T
�Ԧ+%?G��/�j���6f�8�����l�҅���e�ڑ3���V!q�6y� K�N��&�%�Wm�I����/Փ��UН�ג�����l�j]�M[�x�-Y����6Y}k�����m����
q~^��n7b�<�0�P�=�����b�M�m�v�)'Z����ǟ�����#��
g���}���Xo���=����^0V����:묳���F��q����z�i���g��δ|��3A�W_s��m!;w��m�~��jK�uԑ��Uֿ�#�&'���c���3ϼ$�i�4��D�
��&���(�9���:+p���g$ۘ��e�J�m��;Y��8�K����B�u�\<�bEN�	. /􊢢B?n����+!.Q<��]�9���.)��.�v�K�{�@��Hߠ��Cc�:����&r��h"b��'��8�j�J/�^E�v�B�c�{n��R�`��}�Ld&b�I�h���p��R�>+�L� ����\����1���1�
%��d�74ֹlKI�����Fz�9�_�<��3��}��vz���믿.㩧g��mێ�E}������6�I��7��g�w͇�{�L
u�}F��wt�1��Ѫ�=@;�
W&?�{x^���%���ں��U�W�-xw��^�;���L{��'g�<�O9%m�ԩ}Ə�������.[v~aa��c������+�R0��� ��ޔ�s���SO;�Y8�s�)�f]r��iW\����������Cҿ�����~.c޼y�ɨ-�� � �$�������Ѧd��1q��ڞYY�>N$f{a���pǵ���B�����E�	�|�ş����v��Q����,^���?ؘ�@9�&����݁�H��|����~�\�M��������A|�6e�K�@۾��ں���ZzN��L���_[��
m��8KH�$BC9𕐴t��I�P�Q��=���ް�Z;�,��D�2�TyɈ�6��Y�'�R��[�k�[�ڠ�l= SA� ����K���N�	;f�WD��(Ql�ݶe��رK�j�+yO>�������>��(j<���+%�5�v�T9�n`�̒�����3����&����J���Bk�B�zW��_%�V�$���j��4H@vH��5Ƞ�k���ܲ���^o�**,�o��x��acF�<$��`+X5�4Yqn�/͵-��۾-�exs�a��GbĜp�qv�̙^%o߱�y��7�`� ��'q�')p��4e%Su��櫜�Nf ;�[e<�:Rd]��D��������i���e�͒Az�ed1�_dcǍ�|�b�=º�*�--.�7%���+N("�p+�+���w��R*Q������%d��Q�R�R�<�����8\
#w�0�����0,���j���i+� ��qgR�W�{S�V�:�����f)h�(���~JN��� ��Ğ��3fZ]�	Ghk�nf�#�H�܁�*|&���Z��:�;��X	`R�/�cC;}���0�5���'�u���
*㑬:�;�0�qe.,*���HY�WS�o5��ŉ���Bzxh�3�f����P�Q���(��-m�_�ǅ�QNY1C�$${�x3�D�c��G��-�BƏ� �,/��;�cepА��gxIh���;�z�*���@�m�Ecݬ1Nг�o��˻��z_�9/�d���7�̉j7aˉ�|�r{����ӯ�O>ioɐ��e�Βr;c�+߼�2m긁�E�-<���x����
����� ��Ƚ
���&e�ځ�{��gm���k�ػ���y�z�A}�-<`%�9Ɩ���,�oO=�����p��$��fkji��?v�`=Ğ|�i��v�Y�g�~�W���"��uŊ��t�i��+��"���:����=c�j%^���FtE$Ο��gnD|���}gb�������f?���ɧ���S�L��-�� �a�pi��(����R}d�F0R����N��g�
)��	P���S_��%pwap� O)��@�w�}B%���2�&V�*����u��Ê�!�#tJ�ݏ���oY��@;�S��� Ȋ ��#�O���{����?�}hC����|�$�&�l���9脠(��2����I��=�I�1!����Ơ?�X��{�=��z�iooM���ӿ�o�~��?��җ.������GH��9�lB���n��D�(�|�����(G��`��D��t�=�V}��ܳw��M�6M�.|�x��E��x:m�u'�ٳ�t�vz���R�y,�>|�S4�~�t?U����ΐ~}���N\�tѴ͛7��r�w�?����J�6�����|"K�t�U�&IiɌ�)b.�5�!�(�0~ ���D��K����9(e(����a������3 �ۏ/����	��S����;( ����ْ����g�U�ɖ�r0l ������7������C��V��z������]�F��$șݞ~�4��/���VKL+�Τb�WYo�R�[�q)H��.}�ͬ����R�ʨ�=�6�6�ێ��,����o�q5U��-�2M9I9ѲJKm̌6h�K�0�Y�V�f��QaM5;,5)���-�N鮰�CE�B�	�Q�N���	H�>�x	��LI �PdQ*�k���>�A�R4l�(O"]���{��>l�<���;o�mܸ�6�F�i�������IKʈ��*T��S��������MJ��Q#,A�h����&xh
�Ʋb@�bb5f͖��ex�ݸ�v�[.�F{�pG�D���>����6)�>�3EV�"����D��N�D�9"�{�E�AT��kͮ�z��(���
����q#l̘Q���a3&�ر�mʔ�a2r�e��6m�d�eD����/�vꩧ�'?q�͘1ݕ���|2x�nھe�f��&	x�+���6ډ�I �H	:�� W�3a�QJ�#�����q�J0�A�(|���h���[�J��l�33��l��F�^VK���>\^1zc�@����1�r����R�FI}�2g���o��Ҿz��6m��+J�
wEVtvj�1ZQ�Q���I���.,����n��a^>3��#����s��Z)��w�u#�o]IR9dƃr��������VƉ}Y�v��p⮗�a@I�bU8���+,����e4�q��J]����9f��QY��~�o�I\��+�+��S&0&f_L?=f��I��y�}�7m�t�q�Op��@��+Wd ~�L���T��������׭_���@��]�e��Q"|g/���ْ%K�m�UH��0N1*�Cx��~�+ihi�͘4���WZ�:�^P^�y�N��F�uXE�q�>&؀����+��o�f�����a��^�Z4�эa��;��Dw�f�F f���
U��o��۬ �9ڞ~�Y��.W�sr��[����2��������2��v�3>��3݅��;��y8+/��(^�`�|��7d`^s�5~�<��;ﴟ���6u�T_�5r��8�I&��f��Ž�Ȅ���lB"
���)�y���#\j�ez�AϬZ�_P�?&D���Kd�z���p��G�G�!h����b�(��+�)�Ǡ�H�G���z������jQ=��?��s�<����%+�Է��w}����d�4�t�L��1D2�\;#�A�4�|�2[�����`�P�~�1h��Q��ݪ��*��ꫯ�<�����G�8?M���~��̹s���K/����҇q`E;z�1�J��D�(�|��>j9�?�#�(�Ex&�t�#����N~��I�����Ez�$;3�Tx\��Ӆ_�G|O�lV�R6�zp-%++�P27��oI=�'Y�Wru���?��G?���;��@�K���	����̈H���D �x莐!���L�!Nf9�af�!�<$�LP��	\�n�w�q���~��s� >�����8�K@�0��[���8)Q0���Q{f�?��3�|u���E�)�g�����������r9v�t�+.���KL)���4k�����M��6�N�]ʋ�pl�l�VW�U�bsW�%� T��M�Q��
��B�Ǝ�iGϰ��>�eo��WV��?��e����3b����l�����P�!\�T�����VP�3�#��a
'F.ㆁ� �9��������ŎY�#�8\G>��׷�����ޕ�_�����}���%VY�ߣ�ܺ�V��b�6�~ì;��6m�p�0z���0�
K�,G�K/��I�PQ�L��%�/�)k�2x� ��8�N���lq�}��.�4	���z�ڵN��zKԸp�:B�,\e����rv��k�=��?#�x���nH~��d2�x�Q3��g���G��a��PN�N��q6i�>l��).��#�sl���6q�85j��_��V�\�+����=?g��qǝv���m۷{�,w}c������	u1���;o��>��{�Q���?��s]-�{�K!m:�B"A�ٹv�p/���=�Rd\a� �}��Ii���/��4p���Ay�3�J$����Y�Ÿee�gI�r�MZ��}��*�ߑ;�1((�r�H(h�������j*1�0�3�D
�~)>(�Acee�����.�Cʦ/�O�=�0��3�?f��7�����v���cH�Qv�އH�{R���[&�0N�l��e�_����f��i�@�͊�p�"�@Lrp�|�$ m �}D�����2���,&^r��}=:a�e>q2j�p8h@41 ���#���.���j�Oj=���K�P����X�8��_��Wv�Iǻ��k���U�����^|��x�u�%�T��a������ַ_�����⃢���%��'<k|&͵�cX�$_���"�P����3�Ͽ�)�G�ɲCl�ڝv��%2��-M�@�`�%��-�`e�D�&�P�qٌ��v�J VAQ���Eu�'ظ�쩧��muy����o���GE��O<�W�)�)� �X�8묳lĈQ��/m��W5�#|eه��.���/a�z��η��؟x܉�}�Nxk�ڽ�ی�4�ս��+�U��I�h�!t>B�nD	N�+/{TKFvw��� A�\�P��Q��X-���-��%�/��\hj6�3�f��j�P`r���B�,�9ʢ�H��ǉ�Q.�}՗�}�t���<�����;�E އ��AF����>b��7����0�s��$�$�$�KE$S9p�1���`2��<��o�m߉�l߾���+W��t���/_>}���G,^��d�#e�HKόE�#Ki�d,��ik��7}�r>J}��!������70�J�ہ��d6������ŀ�g�PNģ#�o�G�TcW�_������u�8��K4���?�E�k�+��@�K�����A�M����@���PF])�&2�)��7	&@����``�\͕�$��=�o6s��������;���?'�n�U��oC����i)���f�:����0f�B :����6�qt������[�=4�c/��Z��/!w���[�ضݕVU�i5�)��R�#.ɚ$���Ų̪��!�I��T]q��J��:N4� Η�0J�I�aV0����s����6j|�5�v��-��J
s���]�'�l�W��l}�2m��y�ԣؚ+l��56oޛ�ּy2^޵)dRL��#���M�B���g�w��g`���\��Q&D��p��l����"%���xӲ3�l�;���"K�� ���V:f��i��}�����KY��Ͷ���*�ѯ��dpI�,(-u�0���b��-%����.>8n�p��Q��b����N�Q��P´a�f۸�uk8��ۉo<�A
,+�'�|�ʎT%���9p�:�79ЁG9�8���f����>gk׮�(sl��Z�8�0:x��~�ee�K��UM�ֿw�J����{��]�@4�YF�~���4J݄SG�pڪ�s���M��y�����.���� �^�ʟ���oF��%	��o�Dߘ5F���a���#���<�>B��(�(�q�_&Qx��b�#��;�e��;j���#%��$8����.ω �*���W�V��̨�ј9�茔fj1x(/R�P6�����+�6Wcߢ������O��yڎR� �������ٸa�+m�)A�l�}���:�a��X{7T���SpR�b��Oڊq���&Xi�����p�o����sϽ�׿�M
��l6ֻ���2��Ft,Vd0�?J%cB{�eO�L�҆D)ʬ��+	I�2je�&��K���I��b��/Z����^��"�i�#\�Y3v�]��/�
d}C����K���5b���&&*�jFT>ʘ��l?�E�}��[�`��b��m\�0�̺�MKk�ޓq+^��]@2�,W��� �
��U��ܷW�gsȴ�:��!�E��*�$�H�"�Xg�2Y<�f|�iV����fٴ��4vs��=�����0n�9F <��]���>1G��2�vCcĈ�n�oݺ����/~Ѯ��z+�g?��M7���j_���]�VCmŪ�v��.�'ex�����zξ�7^Ӟ�YKMK�aH@�h��'8A�Dp|���l��jY,�}�q(2�謄9����=��7<yh��,V��S� ��>5���[n�����܇��I���~Ԅ)��2D@��o��+լ���K�a����'|����!x��O7�D#��v�3��͎}���3�H]����'t�q&4����R7<�+uQ��B�`�.�f+g�����Y��e�����xD�դ�whO�%9�o�Pχ�׻-����?I��7����qTf��D���_�Y!=CW�P�%�6D���^�`8�(#���~w����>���U��W�ǚ̿��+I��ALd@�D�B���P�|`qf0�G�p�A�@�B�!�Q�P.0��Q�>��B�yR�a������Y�!Z��i�
��7�������v��!��Z@��) 0�P����W�]ӫL$$��`����[ʫ�kc[��]BpNJV,kCbp"i��6S��UcF\M�v)Am�)��1=Ϊ�:l_S�����ζ�l�;+��f��k�g���Q�}LR�U�f�ݏ�e7|�7��칶QJ��}��PQQi�-�?��.������s�@��F��_�
p����6��7	�3&��`4������j�j+-*�~�%q���dmq*OL��;��N�Ό+�i�!�nY>ty��r�(��Zy���4[��I��e�oXe�1���"��0�h���1
� ��8�V��e�X^V��UVٮ-۬K�<-�T��]=��c�D	\e�:Dk�����8�E�4�������o�����~�=��C�l�R۽w��5T$غ��2�b��W�|ݾ����/_fs_~I�R�m��s�	'ڏ�#�<���_|�^|���g>c�jw��?���2h�qwԴt��D+ 0p��o
�G2|�~�"��5d��e���!� \8k���[=t^�?(({D݂�`HQ.����G�KKJm��VV��K
��%I)�9 ��R$�-�z�����KyK��=m��V}P���o�(7(��=����d�.�"�d�������}	t�~,Ȥ*����#@C��Ja� @讎nKKM�a3�W��U�1c�|M�P{#�J
F'J#�l
E����}������� ��Xg��La�K�7	\@�d>j{�:O[�J`Kˇ��Ӝ5�q�s������A��?���3�/�j���7�?S_}�RW��dr��7��7A1!E
g�R��`\����8/<��u8��sÆ/�/W�E�'�@�C>01�Qm�OI�khk�'���_mEF:�p�ou�!�d4�Q���K�Δc���n��f���}�C���B�^V
�,�}po��|��{������'c��y��2��z啶u�f����Ę��j�rD�[��djj��2n]��r(2��hQ��%�=F��E3Y�O+X�x���Sn[d$�]�V�,�$�z�]��N���#Vڡx0�M?�IhZ���YI����<��=��s��J9�A^�=����;dƓ̘�h�rho�uk�ri3m�ʘ3F�����-�
w���G��~�7���ڬ3a�3�㦊��)�6`XR��b��h�y���H�l�f�B�iKȡ�?�[�����?J���'��~��'�d�I�h��E��+��C�%�粡g�)/�*�So�#�w���+�N!,�I��w��I�R���IHHS�N����� )Cf�!̀������P蝩��s�3
	{�8���W_�[o��]����]8�P�})�����ԭ꺨�s�A����)CB��M(	���*�d,p�CS[Kx�3o�\);�R��$�X�hlm��U�m����F�M��WgkVo���Z)��&ypY��<|���o�Vёfk�lGm���[S{�+,��d��^�k���Wc7L��|��x���M�1I��L@�)㏀dƗ ����<+)�c%�%j3gX�XsW��u'�֚kK�c2�꺓����R4�YٹR�)L�MV#c���Y�f��K�WU�8��)�����>��wI�j�I1>��$��Nd>6+'!06�aA��Fp:$f ��{2�=��6E��g�.P��BY����ޱ?���v��7�y��.1_��e����l�����;��n��>s�g��γ�y������u�M�j�Z�����^y�}�k_��y��"/B	ٽ[-�*)f(\Я+�̠�w���� QcJ����v~��G� 8��z�J���� $(Ð�!�,0����GBE��{��:�m#��&:1���IC�"�5��>�&M�P~~����M���VxU�+�)�"�;��D�#1n(��ڎ�wo��kve�p������]�Ĉ�e��<����#<EX���D��ѡ۸�F"�����,��D����8
�����+o���C�։X�JA
��r\q���ٳ���/��]�p+���UUU!�zBF����/p������ߞgK�.�-�7���[mǶͶk�Vۻ{�mX�ږ-Yhׯ��J&e�l�{���_��n��v?����8�W�ix!��Sl�G���E_=�*|?��
GI��CI�=��#�X���?]1�?���LFĳ�%�p�L���C���I��vR���~�Y��Пḧ������}�y6��0N?�+��=�p��p`��'���L$`0����sα3�8��&Ep���8x��������O���N�,�ļ7�t�4z��	N��JH�N<�;�hw��8�ޡ)�(�Ɏ�))i>��D[YY�l�ڿ�v��-���X����m�_��>�z�8'��ܹs��Gy�WgIOF�� _Y�|��ם���G}Ծ��o��.<���n�C�Y=>a"�>�F�L���x���G�Z����h�.����Pc�=�2\�����G;x7L�����w���O��:�'2�9+����z#s1v����G�*��������!ǀ���bR�v�L��}�#�:�?j�]�.�.�jxC!�[�ӊ��(����q%7�~��'��Ɂ6y�GFv�N=;�\�J�z���y�ڵ�&K��@N[0A.�Llƌ>��	��;E�DBf��"�!�wr�0d$	"���q!��`�!����)�o=@�"�'��ϊeD��E@`�	�K�o�.�z~+D>4�=�>�x߿Q�%����CJ:geL�1�j��3�2fY}�+9ݚc�]��~g$�_(-"�&)��~�i�ʉ��A:��p\�Tk��q�Е`ɱb�"^�MNͰ��茕�#�mʑEVYk�����L��Sl5UR�����XK���P�PQ@wI� ���3���p}�yR������yb��R`~( �?�{�u�4٨�#%�,b�0���Y�i��m��,o�T�v��j�-_�T���7.A�EB���)�� �qo�� �&�8�jC����N6�n��1�n�Z|B����[Wۮ��-'�4L�i575��c��s�<"|���]ߗ��a�8�8N�u�
,��1FgZZ���\)0�z�D_�%�W�:A˗��ŋ�آ��]��R\ R.u��#Ö��E����E���}�g��2wa$b�ӞW���`F G��R��ϳ� B@��=i�,x��)��te .�]���"�{�ഌ!0J�3�2|�WY�?2���nt�]n0�[p�:kk�^�5� ��p7:\A�e`O
BE E�p�(�����06P�������>WffQ*�=�(���:�8�Q�Mڑ��'.��"E�}��T���vD�F�~m���#8c0S��M2����E!.�2儲�meDW7r�h#e�Q�9������9Gf�i7����!Z�GIe��'+�O=���O<�o�'H»�.v��(�\6�J�}��9ω?cs^�c/(?��#�|??�Y��_�r��^<xx�?�O���):�V{�?t�9g{Hu�m�x��z��+��+����ڹ��O�臨(�2	:��&:��Sg���n��Xk�F�ۨ�%�~ǡ�]2f�@� /j�2��%2^�E&�;�����Za�-\ku�1���4K�+�t��^6_��bm�ɞ"𫺊���EԵ6w�;��e�-���n�(�'N����ڍ#����_����
|��� �<��l��{�.7:�S�I'�hg�τK��a!��d��Wʝ�iL�F�`RY���F���cF��g�nbl��E��+/��4Vz�3p �����l�2�<�\=j��cIi�d*&���)v��'��5&28R�w�h���2��=�˧L&�x#�� IFA��=+����(XS�B��&��?K�9eB��M�*{�G��H}饗<�
��Y�3�	�
߅��>���y�{$x"A���h��H�ݢᥢ�%>���K����t���&*��6�?�t�90+F��	�N�o� t)�=��+&�2m��7��R�g.��;�[�d�#����V��C۽�!�Ük�!��y�+����b_CIq��3�8c��~��FyR�ׄ����R��������8]Ĉ�	�.��g�Q�G���$�
�E��
��E�q�9��yA@�+��fk�M9$)j`i^.�SOY��CӇ��MO�� !L�cr�Y!�dP_e�`�����l9/$*��J� f.��E`'�$X���u�N�1'e"S�;MC�U�6��#����1�o��m��(�5l��֝6��WǊa��L	3�5Օ�P_k�����i��[fk֮�8� ��+3���(R{��6E.=.p�*,aH1
�[��퓠.�S`�2�X���O���L�o��}��S2�J�N�R�V�[&g/���i�KQ� P�*�#}�[̛��;Z�[��s���J4��!I�.1&2 �D��jS9&/cwN�#�;(�$�I���$�x�<�xۙ&è�!��u�A���?8���U6���q������^�����II��u�`A���6�Kyᛜ�<g���^�2a���9���}"�� �q |ecq�\ C#Z>�;h���I�{�{�	�A�0�#�ˉ�[���"�h����2�=�n�D�{L�B�+�g`���Ma�|劕����a���Ir��ۙ1����l�02���8���;�ð�Hcf��u����;�Ĉ|Fhv2�E+W�rc��h;x���(3��O&$6
��S�N�iӦ�L)���t�ev�����-JW`N����'�p�q9����'�ё��A] �%	ܡ��CD1&K��F_��翸������*=�УR_\������A���(_�}Æ�2^V��:���m�D@��>V�7o�Հ5kV�B~�̣?�e��}��1S. :�Ga	ő�P0��æO���z�}�/y��AR�I+W���v��G�'g϶�?�jk�̺,Qpr�	v�8I}L荈��x�t��1����>�;�4�t�m��`B ��{�|�;ᤓ�gD)2���$�bX^~���{Vi�0�n��!��F�0��.�s�=v�m��!����*��%\�O�N�����:8���m���~2rƌe���7|��w��ch95%��.�)����&G�d=��[���s������[��sd	�
z�d��]&Q�\ꮺ�*��/~�vL�4��t�*�q����s��.n�;����H����v���y _{�
�	<&�G�>j�?�f�CC(�v$�c-]}�3�NC�A�7�w��"3#��H�M��$2ޢ���������>�x!��Ѿp?�om�h�z�?�	��$74�QW��SV1��0�O��+�W�Z
r'��J
r,����D}� Ӑ�k��#������}&����up���I����&Z�P ��z���,�G1 �'�L��	�	�e�B�D0���g�	`�0lR$�Y�F�`X�|�bɎ, ���9$�$9Sgc'3�l�%
PJ��)�H�tK	;�q��SS���I!��օ�r,�"�0V���e_c��9'�ߺr�]��'�>,Ѣ$e�fXN���PG���d�+�����$YR\�թMUbr���ԇxQj��b�5�j�M�2�"Bd�\poj�}�Ю�ʉ֒�g�m	���f�]��8��)�o��~	�;wX��22�d�^�k���d�e[{k��5��6T
-��o[*��;�Z�yBhwjl`��-�r�|��Eo�2��9Ψ0���d����[Ƒ}#�����-a'#WJnCw��L���V��h��T]�wڥ�tXqN�..�)w�]���luq-�$c�#.R`Q\nk�x����$�L��8�0&��q���?1��*X5"��hҩ~u	-��.60��X��1���^��H�6p�w09M@�$��iK{G��Z)�����ڭ-R�k�V�n^l~���tc������+T<��D�A�z)�2I������xQ�zP��*� ����p3�&0��=1Q�uO�'nv�!���m�H`���gQF��INL�MV�P!C����mm����P�(v��m�mR�P�:�.U�zc��tk\�8o������{�X�}��Z(^����*嬡����J���x���6J����D{0�4�R �9�]�+WD|۸����t�n۷��u�x�J)��l۶h����-�E�� f�q�?a��<I
��Cm����o����6`P����+���)M1(��T��E8�����!�#��0��1�1�8�X%o�;�x7n�G+t�P;9����7{�AE���.W�R�>��UZ�O�P�ce�YII��y�}�Oq?�W6H�� +(,Q��� �}��i2v��g�e�l�v��h�O8��M��ݻw�؏V~�e<��_m��~��v���?�~�����'� +�բ�oH�߼y�]s�W�$)��̜i���3z;E��%�ZZY�o�3�:cK������T�6պR�#>S8��V�����n�;q�U��+T	j��部�������SNu�������r����	���T�����f�<�F�k_��W�#g�}VNp��B��"�Z��(	Y��A�O^�I۰~��x����=�ó�<g[�l�ܜ�O�#��Z��Y/���~�A+V/êc���~�j[0��Q��'m��]�i�[�q�m�.����֪�����2�<�5+X�<�=�������|�o��S�۳�?k.�5����իmي����ٝ?�͞}�i[�d�-Z�P�
#��ƍD�j�{�-���E�WĪ�7	Є����{�.z��oXc{��mn��N����	޼�#":���{��o�rDw���d�ƚ�x1��a����B�;��8����eR���Aَ}�A��ஜ"=a@Y?+�ͱzν���,j���:k���&ޓN�(��&}H�t�v�
�8������N�6&�1�:d ��$c֮,�8��z�Z۸a�~o�%����x}�`�<������"�S0 B�?�����)+��+���A
|��x'���?�H2���	�LC'����	d}�G?F�oB�Gg�9��/�M����h�N�2�뾞�q���;v�8z�ƍ��̲����"�f(N�33�:���ę!���\��%a'��7�
e��������3��i��=3!,�v��.�������I1pf qMa�/
������(�~2��s��L[}vV�MF���k(�D��=�cfIi+�V���g�<]"�Xe1[�l���h�����ʦ~��!��B�o�W��[ڰ`�.�����0�ӦN*��<1�*[�d�(? �E�@}�%��#���3��6X���D��3�EI|ª�<1���'Z��2YF��wIx-�}IR�o��w���t��c�;ޕ�65oպ�.�2��-=+_�\�յ�۶�&�N�c��ni��VQ[g�2��e��W$q��|�MN�j*o�8)d	j#�ve��Z�O���gрE���P�{��Xc�n��r�f�*ý =�v�Yj{7�g�f��L�=M�u6l�p;������Y$X���w?d6\��H���I�p�(������w7���5k\�"p�R>��-Cƞ�c\
锏���=�1�('d)�W�ۍC�*}�xM�|��p��0m\p`��#}����G�{x,��e
�m�����H.r�����q���-ơ��mzU>�О0�L;�y�$wfnq�ň�~6�'�=,��m�a�(#:�^Qq�53l�I��� ���:|�F�
�bbC�Wq�&�X�a���W�wh�4!$�����/��s�^6ɳɚ{�+���C�w�8E��D��%�N�06]R��/��MT%Ƒՠ6;���=�{;��y�J��8�m���ll�	'Θ4�QW����e"��++P��C���4��v����b5�`
�\s� ߰B�{��؄:Q2�3�a�\e����G~�A�>���,)%���V�vJ��|o�k��,�ɰ�/��q8+i�֝�28x`?���t�7]����Cl����,Z��H�jGl�5��*c?&1��3�M
j��P�މMJ���l	)��[�m����2�m�,R���γ��Gy�L,�a��g��J��O_b�������k󬶮R��hU=���{q�|�-����������9ϯL*���裏�1��-<"p����ƭ[����q��6}����J�~����G�W^}Ş�������<p���+/̙��8�v���O<a>��G d臷�f^t����Ȭ�77� 2.q��n��7h�lټ��q�ŏ+��ĪZ��
(��j�� �iÆ2���bX�׬�}��-_��`����)7*+�O+*��d/� �:���Sv�z~��L�����I�Jhq�Afg��j80��Xʧ�Ag@~��{F���l�=f�h;���݋"����:33ͣ@�vr�Uh\b򙈝��r�kt&V�X�d�Ĉ#�t��h�i�6v��>��3��:z��O<i�ԩӚ�B�����F�Ӈ�H��	����9�\��A�4�.�CtJ�����O&�,����\�|KY��;�F��Zt�ک�����;�0�@����O:<��_z�+�n�Z�aD�+��ނ@�n:(,1c ���a	�@A0�@P<(��d������j�F�������S����ކY���>b��0|�ӗZ�����w��{BY?$����NoD�@rfv0��(�ÿӽ��x�s��Ϭ�u�m߻Ŏ9�4���7m�>)X9���hRJ�-��So�Z��q<Ӎj��KJ��k�èL:��1�de�
�ӥ�īY2�,}[��fGLͷ��[2�����v��'�o������x>b�M>�־8�����'�XQV���[F����v��h�O��>�y�'�c��'?�������77'�ǟ�r�Swg��ݽMB9�n��wm��3����^y�M�ͯ~ci	RP���*	��2�R�l���,6���׶Z�|K��5)-�ʖA5|�P�--�v)p����]FY�2�#{��
3ZL��Kq��]�tU��r�S�]�S�{�Ơ]R~V��O��w��m{�ˌ����&�L)2���9�|��?�V�/ԯ���Uc�x<6���/�*��<C����㏷��Ǻ�
� ��H��L�ڵӅo�� ���3eD�Sl�'��FC�:�ܧ�	�T7���X�봏���~M5�w	��9�)���e�1FϽ�/~zs����h���t�WVjY�����%5�7t(�#V0"גn�!�Mt�m۶�K-� �:�F���m�?a� �E7���-���-$lw���U�y3D����	*�?�	�73"�11�B�p�"w�t�Ï�"���<����~�D/����
���Xp�	#�p��s��a6h�P72؜N��+��A�k'p�Ɯ�`V���N�᡿���<R��w�]y�W��Nsދ�cЇV�0��My��{��rϣ��h�A��}~�8���Xqe�ͳ�K�����NINs�B��^�COW� �0�	p���U���^�����-�)�����,o^n�=��v����G�c�|�Sֿ_�e�'��*�묷sO=Ǝ�5��j��Vn-���d�oh��c֘��g�Ӭ<	L�	 ��g�M5��l�����~[�e'L��t�]vɥ�Zɠ�8�~��]F2�=��:�����E]b˖Ϸ�*0dOZ��o٭�~_������j_�Uɐp�f��p�X��5W�m��Ѝ��|�
�?���?�k��A_�U���~�*{��� o�-��q~�*:�>d	�{(�B9ǟ�R��1���WI�{І����䆰�{�}�AW�O9�4/#*���wVf�ӧ����c��M� 7���5��DeKs���L�\��2�F;�wʋ��;���,�tTW��D����K�x	>񭛿-���ɲe�y[XA&�^ԗ�8�s�z��{]�Ox��W�f�>h+��7���Ǌ�c�ㅉ-d{�"��t��p��f�QȂ���Z��k�c/+רE4�Y%���.[��g~���/����N�Ȃ@�!u	6Q�&��_9��K�3��7�	-���y��L�����3��f<���l2�2)\�lV׮]�u֬Y���W�z(77��/qO�����t�ץ���+�͝;w��F:�A�$��� E��a3�
A!�QPP��e��>���
�#��`N1�����rf��%{���|��c|��ef�~R�':$��j�.e��C����z�y�ߞ��z�M�}�h�F�g�����"�:��>H�Z�~��o�Ⳮ56�:�Uf�\��%&��Be^zyT�#F#U3��%���Q�����.�4&�FȲd������+s�Z�nGRY="\n�h��r	�f)�����ج��%d�T_���4wIk�"3Tm8v��-3W���H�"�کlLg�F�&��xH55�:C�q�a����^�ƞ�նmo�մ&ٞZ1��'k�ye�����+�|v�[�C���dd2��QQ~��gYj|��(wJ���(���GN7� eY͊���\����ੱv�X���Ȕq�n�kָ{���Kx#7�-~�i�6}��qƙ�cĲ�J��G�3=p\�iWP I��9z�1v��a�F8����0`�T���8˗�WP��ݗbe��w�)&��{G�ک�e0",�MxɌb2��;g�o�)�מ�0��6!dQ�[$�Y�����@����#��L�C�Q���C��4����焈N�eR�Q��-�0A�:�̔�tf3��L�x��Y���V���"��*2�÷r���q1[�X�gFUU�J8�.ѕGl�r���1���L�8I=�q�Utxe�Ǹ��@�'�IF�D9����h_"p��%pb�� Q��O�R\R�3��<�F�_��<��Y\(��6�9���|���p9b�1jh���/8�&������\7x}hW�89Z���
=0��c�1i��/|�~��zd5����c�SYm�q�F�F9u`���~�9%³w`�_P��
>3Q���T��Q<4x����/���,R�׭��+H�u�N?��2E#��֮8�SYkM��6v�Q6l�>�3���l�8k�ť���Q㭰�P�((��¾֕�au���E��x{o��Sq������϶Q��z�5�U2@p��DѾ�B����?�W^a=��y����7��;l����n^G��/�(`��MV�N��n}��P.���9H+W�����=唓l���i���=��s�j�
_� �B��"�G���J"����Ô�{�!VS���h�ĿD dh�e�;]1��f�U�l��t�Y{�X�ԍ{`dl�9h���y���9�8``�~�br��Y�G�@D�u�L۶}�=��3����=� ��>9W�����3�Z��p�����ފ���|�~H���LF`Ȇc�n��<��P������f�HU*�Pd���*ωڷC��7�j`Xa��{���J?8��7�x�p�G����S���>�t?̆uk���O�?�����D�I{�� BBG��-���~�~�o2�	~ �;r�,��|ލp5Za�8�Òo»�x�"9ώc�^U����'�|�;���V�W�w�I�X!D���Ddpr�AFh"�D\9hE�L���Of�� �A�U��H�@���!Yz�`�()۷�Øoo���-]�Ė.Y�eL#Q)�+)���3@�������;� �F���͸RS.���MWv�X3Δ�s��}j���X����+�<Q1��#\$t/Q���L䵵K�����3l��tk����_ߴ��o�;+eH�<��NnQ;��m�aGXrv��f�-�^n��m����e�,����i���m�)�_�P4z�������S�rjb�%�I����(�O�S�}�C
��Q�۔K%Ц�<ޚ
l�iţl�̏�e�٪m�VQ]o�R'u�M�5Ӳ$x;+�-�U
c}�m^�Ɩ�_dջʭon��HiL8w�5�n��_ ؂$�G���͐1��,({�P(�h���	�����AFHG�G~K|%A#���A�(�/j��KL�wQJ�������`?���(�(�(>Z�:u�]��ӟ�����O�'?��}����qS,#=�f�+�mMU�U����Z	�D6d�<Tm$�w�5��w�Y`h���Nh�$�zػO!��A�'�A
}��F����g���mǎ�%�����U�VK�o��X�+���ر�V�\��{8G��1���	nrMML��o�NM�P�R\d�o߱�v�-���&���N)��_1R��tro��%�#���#fO|�@�À��� tM�ۡ��	es�`�3���h�$GnR��^�Z����\�)�C�8�I���S���Q}�D4>�R�Yƻ��Y��A9c�٣�)�Q�h�2�9�%0C!�ރ>h����<�7ߣ��y�~��� ����~���yj6���9���U���O;�7�<Dc�@�'�����qMD��L���U(�gi�r��Qw�^��F�G!Q>��3V���SX�ߖ��b�\o�e�g�x��*�
;���V6f���1���JG��aS��)Ǟb3O;�N��v�eW�Y����!Wk-��*E?9-ɲ�{jff4ƣ�o����}V(P��Q�0x�S�YGD�֬^z饾ڀa��/�3c��O��v�ş����|��{g�U�!��uy����*&�,4��2��+%x
-b<�~�a�5�[*��葡ܡ��{!�T�t�2�O���Q��~c8��h͚U�����2?"�d'��v��"�I���o5����m�X�Io�d!
l�Z�;�/~3����X��~L4E�G#�)�		24�7���GK?�>��D�ڐ�����{�^ɖݾ�h�x(QC1���~��J��:S��kW��%&c�vHY? +^t��G`��3���K:(�3�r͇>?4�~���?*�����x��Ø��x�oƈ�<�~��H�\�u��B9�: 	�Ѓ{1�����w\� ��w��H7}��7�x�X1��6I�B�H�0�2��e���;���$ e 0�Ҝp�I�Q#��Aɤ\�F��,��OU�g6�hk<���YSS邐�,�Z��� 1+����a�D[�����=)��;ˌ��7��}�+3B*�[$DR$��0ܷ�@[�v��ol2�Y��v1G�����-�>SvwF� �N?);zO�aH��Ip	���n��1P	��7�+O�n�l��6�-!]ʞ�/�?g� +6���,MB�M�D�\·5��b#F����t۽k���6t�h;N�OM����F@)��5�j�:+�/U�R�E��1I�~��)�jۄiGZ^� [�y�m�Ua�mIVѕo��GZ���VgI�eo��h���s���A6b�6�D4�vo�nR��w��ڊָ�O�}g��.�Dx���#`��3�>(Y�A�;@z�3�GQ���G�e��Rl󒷬n�fKM@��B.���[��Ga��r��A���|�^yy�%I�E��t����9�?����"�r󥬠��� P ��͕1H���)�RZ�m��
�,*TH��>��6l�p��-��n'�}�������хr��a)�dm�8��o�\,���7���dR��#�"���?R�~��W|�Qx��l0
7�:����z�����ľ�27hd$�,s^
�q��{���Ï�������)&D��V�0Ș��(mm�{F�'��6F+pѾ�?~GJ!�/���_�>r�m"��Ñ�Gc�"zM�E�{E��i���@�5��'��
�^�/|�}2�6���>����R��\c�`�2�̞�?���pf�[�m��fq��mJW�_F)g��xf��iӦy0�0p�!�Q�9�4��s�3}��A�x%���a?�2�n�͊^�p�b<�ݳ@}���/�%Ro�"�t�H�����-\��s������߰���ݷ��Ơۚ�C}JJ�3δ�N;�����V����[����Zڻm�捶y�V۲}��߸ٶ��m[d�3~qRX��K���/��2�TWJn�.g��uӞ����sxy�EVH�Զ~XFl��A����e�C�3�ط3|�H7v����aU�+	X��|�A���o9Ό=ʞ�9~�Eڐ!��}�g�yN��
�<GG����w�`�c2�R	|cܐ�Ļ������[�l�r���s����c�,�w���x?-��䓳�׿��m޴�W��/�@;�e|����{��H$I�v��":o�<we�e��%p��5+5N�m���p~�ź��$���˖�W�m��A[�>��o��I�I{X��
]�~c��wޙ��
����u2�v:�1z�Y���:O�&Q"�Nw��̞>��t�=���?|�Ƅ��\��'h��?��l�82�q���m�w�c�}�F�MI_����W_}��{�-.)I�I�+m��2���'{>�I����}��B����GI���}X��GI�7���5��p|��Ox��Ɛ�wė$/|B/�dG8tG�J����+++{��SO]q�wF�+��@�K7���1��/^<VD�ᵈP}' D�$����@��g ��,�"1��� ��eF9"��7墼��ddd��Ł}.`�>�7����y�61�ˡ<�:B]!���aO��}0E+G�	�; 9���0f��?v�H���kK�cmq�2����~���jYM銅Y3���P���U���j�,39�vm�m�g�n��*$��%`\��3�$�Y��2���Z��������
��tɨ�¨�J��l��2����U���.�Ys���KNϷ�嵶s�̛�<�'��!�g2�Z��CFTg��rV۲��^���Vo�"�g��Z��#�F��(%�EJzja���c��R战D�-���J!me&N�����p۹~�5J���ϳf�C��+x74N�S��=�ٷ'�CQ|��"��z2��@jػŒ㤐��#�`�-M>�z����fWƙ��[o۫�̵��H���0�ѝ��"��� ��ot�駻���+}����h�%�gRW�"�^��B�-�%�ߓ L�}��f���=��9�\P6�.��B?�d���>�芘�iK�'E����F��)�Mfs��QڬnFF+$���ݐh?J���Q�m�q�  �wH���o��� ����ԅ �7�O�N�V�"���t���3��~h�ǴU�f�b\[TN,�2'E�(0��3��B��� ���a�A����0~���4�z��D9��$�� <x�3�KX��½H�d5
�K`�	�O$�i;0!���=���Ճ����v�;�ڼ|�27�9'��p���7�,V�1�H�`e��b1rx���B�c���s������j��U��r/�=Pܣ����HA~�݅V�g���-� ���O�7�wx�˲�Ш��!�-��}	����R.[�^a �9HO<�������6�_v��v�ş���\KW
ػ1x��E�%�2A�8�(��Jπ�Q��I���o��+�eu2N�<y�'γA��k�j�nW��dC1��q�{Tmk���9B��c����D�0l���M0��E�����v_%��_�z�{u���!�%%Qݻv�{��v��U���CD�Ę��L���᷺���i�)�κW���+|��駟���_{̓;̛��J���+s����/)s6�M�vlM&��j&����8>q�FF>+U�g��Hv��R!���f2`�KsՆg�g���^|I��l�׭�Iԑ�Fy� �7��i����3���g�͐�Ϟ>�-��b���F��%�p�	��z������D&;�`�\5ƒ>�{�zVT�.u�k�&�c��ǭ�w���{/�O�rrr�|��3������ӫ�����X�#֯_?���$�1����8����C�z��;������g����)��;����2C�w{��;d�3���G�`]\O�J�T�@�e��Y�gő@[��������G��@:��ݓ������^��#>.&��Ɂ�	H"���x����/�or�:q�'2��[�4�4~H򶹢�A���dR�̽�>���O1��yT?L?s2ߴ�K	�6�ӕx"��{>��K�dO�<��)��$Z[���o�$x[�%Ƥ[Rr�&2˲L)2#�N��c��x��zBW��j)FDj�-ȱ��Y~Q�5��n�����p�u��V��Ǟ[�����{g�=2o���鲺�b[S�n+v5���V[�����j��{ۭ�!ժ:r셅RB歵�]�G�g�*K��-�QH��D�3���-���,�I���!�BH�QS����-���b$ܻ��]4X�Ui��w��y��g�u�@�d �,x3>1��?�s\q�W��*�	�4��4@�av6�������;y�KR$�"�����(��V����L ��6y��k[��i���Zw;۰q�j����R�r-?������1�FK1Ym���A�E�"%��
�����3gp��я~lg�}��M�����?�mO=���,_s���^�Y�B�J�#x���^���5&=�@4��wcF��C�>�CډVud��93�C���E���3����)f�J��c-ir��KP]��	2�p[�_2���ޅ������D\P�PE�\(�a�-�0�Sf�=������>;���#��3!Bz��>G3��7�3�:��r�oWp�6���,�7\��ff��%�|�g�o��&���o�o}�f���j���o��G�f��p�\p��C)gu�{<'����7��ubTb�'?���7"�r�-v��W�wW_}�}��s���^{��wI�&M�>�W�0�(�x���I��E��Ф���8ʕqx��!����l��g�����X��TE�ٖ��e����qcl�6u�T;����i�ٌ�3lʄɺ?����()h�%}��622ceTy���D_�ޮ�=(N'��*�i?c�^�ǌ��<��jV���߸���_fee�<@����|f��<x�@ߤ�*Qdq�����B��8��d�?&��wɎk��_W�%>�i�Fߏt���׿��]��/En��G&���"ޅjo�2W�Y����h��k�/�*F:9�U��w\��Z g�V��ɬ�_��z�}㦛m���JDv��z��@?%�*c��E��IV�0���^)��5�ߧ�d�,ԇ���+=��7/�ߴ'�0W`N�i/ψ�	�r>��	�g�uX�nnnU�ْ)e�#ё����'�A������G������
�c\[R���N���?��'�&��a���w��y�k�{R��e}���L�[��S�9��o�cJ�ɐ�}R|h�������Zbl1��0HH0f�;ol�,�u�@��"��>��������GH�Kez+��ޑ��Չ�X=󟎔���Q���G������{���e��SR�������rrj�3}��ma�>���%�C�����mT�K=���>0���nH-Mݖ��cæ���!�,�0�KY�r�t+�������p�>����]'�)ʗph��v��ɖ��`kw��&)����\<���
mUE���f�mi���1�-k�4˝x�M�e9��7|���i�����)'X��)�X8̒
�XCL���=u�V�����e}m؈!���*���:Pi�D)�m��6�7l�y��6|�TKL�"����ʬ�����: ��_�Jƞ�a���A�xL�����Q���~��x\f\���k�2�(6^�(=���]�.�;
Onn���jĆ���Rwo�VH0جL�jU\�o	��!�>f	��G��R�̣��D���Ck��~�wQA�2{Jf�tqI���R��y?�u4�+Ǻ��V�B���p��%�"�#�<�����{��C�����fNs�f�|�\ߠH0��~����@��1>�����'��õx�I	A	{ϼ�^������`q�	\=T{�D��~����J�o��~�L�P���%��V��=��M�c���a;�9������z%�
.�b��k_�/|�2�.�3��������.pGy��W�/(�(��(���=����&p��0C����oW^y��y�������~���y�cIa�3V)���(��	?�@mf+(�7�t����pWG��xF3ᑂqhr�C�䴥�;�8�9|�9�	xi�}�g�8��?�|�T�=��3��Ks�TW�`��\����v��l�V�d)���Վc���Հh\0��~�y_q&��#��7�9|K���{���q�Ot���С��pK��qȐ�2F�|�	��t���Z'�kB��/��a�F{�W��H�)K�UTX�8�A�]2�;�$����	�^�a��{h��ӗ^��?�y����wZz��E�Dp]�V����/�rFd@X`A��x�O�hLss�܍#���qI���,�*��� �p��Mߴ~������+�;�w�]�}�����K�%}���J~3钟E$�8�f\�+б��2|ɟi�8�C�}�G/b�]��Ɲ��/5%]�D<
>�D�>f�4"B�!��hà�]���,�?H�i��}+��KZO��2�"7?�
��NI�a�a�|�w�g)��OЭ�C<J�����g��=c�����1�&s�g��C����X�O���@�<��I��i�t�=��V��!�C���=�x��|�p4�b�B�	f�
�B�d��g�O�h^	�6,�l��� J���o�����#�Ą�/��W�Z�*u��_	q1R�#�$�wPp�e%%%M�"�r��5KH��ptxZ�~��l���K�i3
2�d��!�����xS\��d1��_�D+�G�s�atX��ѩo��$�;clE��5��8K`�Ĝ��'�I��_�[�0�;ْ�E���	*�SR�`,P�v
f�G|b��tV[�5Z��6��m�I��������m5�b�Uj�`�*�vH�V��X	ǌ41�T�GS��H�s��m�m��V��h����ކtkN�o���1�q�M��6��W��W]i/���;�\+�u�eL8ޚrGZM|��vd�νM�kO������:)���m����w�`�dM¡��N?3)^�h�tH��2��m��n��>ܲ�h�cG�e�Y��ؼo��������&��ة����6���|1��x�_�`� ��a��.\x/����Y�Ǳ A@���Jc�_�7�0:�1%J�p�~9ct����A��x�f咥�`�74��� �D8�i�{+l��}R��m@��R\$�E[-����|��l��n�v�i���QS$����UJf_���0�ʃx�UU��ӳ���>%eF=�າ�|��\�Զ��`�lW��')��r�y֊"�*��	N
I�Y�ֳ�=_�<�Q�6,��,�	�K������3���1��-��)�;�1���.��D�519R$f@R�e&R��������1[���5����[�A)U1���B���v��h������!���Z2U��T��32�BV�՗8����ظD��.���D��T.��M��Ge��/ �@/�茓Dj�c�dp�`#o�.<P�������� 8���?��^�;l��VR����{=:ls�����HzL���~�:w�#Z�k��a��~{�ŗ����հx�S��
��,=�Кb,)>Ǌ�Z^v?X6���w8g�5H�����[�R��Ed�k%2�X9g�?0�1$e%(,���ç�s�28�g���=��2�[G[��ig�a3�;Ί��l��M��_�����o��'��o�f�W-�����M�&�Q�+pd\c0�d��+ٍ�ӃY��-֮��=1��mQ{#�(:�5J~(���� (O����*����SOًs^���-�s�s��ٞ?�[��ܻ�[�Ү��F{��'�ـ�?8	��gS�L��>&q�/NG4Ε�C��D�Q=��*��m�����OW�E�*�=�ݽ0�5e�*��������b���)��C��w���a�-��,�����Y�&w��	�E�KKq��Ԁ-��V���'X @ �ͺ���>sg��ʷ����9��}�yFϜ92Z̀"��d�ڬ�V��NeI��,[��Z�j�U��� m=��u2nk�V�WW)�h`�5V��2��0[i�J����`���z]���"��;��%�}�p��W���m���t~�i����ɓdx?nUUe|�)�J����.�%��}�[]M��>0�!��ƞ!f��}��S�k%+��f�*��:���,UY8A�Ix]dc?��&O�,�/��W~AfsAa~�� +#�IQssk�-���a�B�����n��~������G�-�:��E���?��ЯI��o���O���K��!�j�SNq�B�c��8_����;���K�& �{E�l��dFu(Ke���+�"��;&	��off���4.Vw͂��9͙��p������bR���A�+�m�[�����@'�X�hjjN����iinIg�Cŵ0�� � C�@@���! )�޹�#x&.�& �B�Y�)u	�KX3��#�RP��0c�UE#=��ev�0;!y�� #[�#/��Qh�c� ���0�<{�$�) �0�NG�����xx��7w���4�q�
�%U.��C$��(r��l)���� `�ʓ}6,��h�V�o�2�,S�R��V1�vF�
�l� ����²
������,��o&O��sڢ���D���S'I��G�Ο7G��R�o%�zZ79(0�6��_n���9߮6��0QF���Y�f{���ڪ֣gO���̀/�$��Hx�0�i.�g$��sZQ{�'%hV�I��<�xcF���5� >m�D��a�]�b	{7�ogذ�*O�a(M6E�[zV�E���^b�J�w��������S�Zf�r����E����ŋ�63"ˈ*
L����P'a��*�Kl������s|�����;�:��e]���=������$�!N�Ӂ$+�e��ޖI�C����	��5K��>: �� �1��[�5�w�'��X����2:�%������;#��N�{L#�!�Q>�3sC��0s���9�AF���ά�7�|�����b�!��ƈ8{��K����mĈᾏ�p��13�%Ő�/3c�0��Ǧf8�~��?��,5%��kT�C��F.�W*~p���x�����x���'����K/
o�h���a��TrX����n���cie�1;��l��'���}1Ά�3p�I���Od��O�A�W��~B���<K
8������S?�a���ٷO_����@[�upG*@͑z*���)+iq;<:X�3��nB�dvpzW�*|�#�)3������W�4C��wL�_��8-(��R,�c���(� )��a�$����g�T'�
�F�`�&i��0|���b o0����6�hn�B����s��T7�0pI�����ر>�J��&L�_h�wD�GZsdlQVe+--�W_�QI��tF�Uaf�Zep�x���s�C��|�ɒ]엄�=i���M���|+�?i��ڃp@�Nz8����ft�I��N�B9����fH���~�`�2�Od?��%2teȲO��Ӊy�7b������{�~���@�_ )��-��Y�
iL�s#�a�>0���ȓKDa��/� ���иH�8�Q0ah0����ąȈ�@��Q~� �2;'˦IY�x�b_��Sl��I��ΦL�(�2]�9ۗ6͜1�&O��o�<Yi�t�ڽ{�Rk��b2̶��J�T+�d�͛3��ΞesfͰ����b1��3���zO%lg#l�D�2��1�r���Yj�B��S�Y4F����`4$G -�je�,P�]*!R�Pgu��Jڍ"��֋��p��n��Cs]�͛6�Zj�Zz��JqKJ���o;�j;�~םm�v�uFoe#�\Ǌ{���L�.���M�/'�3g+�z��˱��b���~Æ�ЕFٺm`��(�C_��%���vi�b����J�����ٴ�/��A�~�H��R̈!�L�:��T5�@�q:RXW�q	 ?�'\�
~�Ĥ�d�=OL������ C�OS�����(@�;�iF ���Sf�k�a�0TN��k�=$��%�+48tW�	�I�U�6+*ȱ�nw_�~Ui%z��I�u�[��c�e���[�[lfn��W^VU~��	�o�͆v�̖���	A���'c���*�\p�*�Fp�
��'��؟��{���K��m�KӋ~�0*3�G(�-*G���{��#l|�w���;.�'M��x�\(7��i����HN+�E 8M��_r���A������~@,@�{p�P�Y�	�EAα�(��a� ��(w�H7z�h78F�{���������VYu[}��l��״Q+�t���z�-m���Ok���tгgw��e�(�����N�9��}�c�aN(����%: �[|_�ͽ��|�'�xrj��w�-�q����v⩧��<�/Ys�ulȐa��mа�~�uT��1i�Ĳ1��f�ml����a�'V4ĥ;b;���C�@��W�haPB����f��� �5��F����V�y��QB���2.�g~�K�c|�6a	0�����Uf������pX	h�%�yOS���E�`$�.ˈ�u*d(���;�,?���&�F�ĥ� ��pnV�񎦲���L-�2q_�q�q���w�%w�]q�v�	'�Ga�s�����O�R8(e�=���C9�O��or�϶�m�Ϝ��Z���\���gW]u��7�rTV.����{��u���3�$(//��^W�^�o��ZFc��	����D�S/h��&P�ap��зI�E�<������������ܦħ\�a������?}��t�N|~�Kz�'���KFWHסo������%Nd�݌�R~�#���H�Ѭ���deed�h��vF��Y1�SSS-�f�p40��u�r��i|�*��"�A���Ժ�8�4G�ӽg���G�=KG觍m�㎶ïv�������W�f��m��>��]
%2xv�yW�y�]m�-������q�p�|�Q��6���5�j�kl���6_��M��~�O�b�-��C;\��b����u����[��cs�o���N��Je�	È�x���8Ձ�Xt;/	^��8��{�峫F��֋r���eԌ ��2�zĥ����AXڒKl�wm)G)���a�e��[�Ԧ�[hKjꬰ������ZkYE����0�M�,A!%�߰!���M�}�;d��Y��ڜE�Mm��qhk#��ދ1re(
rܣ$V�I�.��t�:	�:�c���o���#ц�KaI7M8A��O���"�m�ĝ>�F���U2ŧr��lF���W���`�zG�c$�YF5�4H~���8�
�o�����O?i���������l��ɶx�")�ٶ���^{�j�쵳m�冢�2:����v�Q�[���|�稑Cm'���)x�ٴ铍�C**�m�_�$!�����3���~�{Nz�1�K�w&q���_}�6@�	�2�UW@��Q���d@��Ca"_������Ge&��w�A�;~�E:��o��H�x&Ll'�����#LB�%�&��a��p�;���4�j�w�o��y���p���o��%e���p�1�͙A��_��W���C=�P����eD��� o����>��%%n7)l[�k`�����W����8 ��M,O���|[�`��hNv�}7o;����� ��G}��!:����Xo�����
��Jr���Iy��r1�2c�T?����F���m���6p�P?V�M
a�8�B�0�I��(�M��K�_�FE�l��C�U�FP�P��xbp���O���s�%��6�e�-i%� (���P�_�N�����D�#�&��E��mR]2�
nQB9��3@UU�t���,rb����5�@L�F�,ˢL�?28�l�~?H�C��b�m85`0��U�%�@f)�Zk�e\S�)<��E���&�n"��w~�ɉ'�d���v�)2t�h��~���A'��]v�%v�e�ص�^m�_��Iv��٥�^j�����OV_���%c��f�G;�r=I�[�}��]����|y��@�Q[QQ���Հ}cl]���������YN�oŶ �]�HQ��>��Ѵ#�	�s���Pʇ�1=��[����0�|0�a�2����?	P�e�e�hc�N|�v�w^��_�z���n�h�]w^���^��_�h����#r~cc������}��҃VH�$���y�>�E�oS�~�@Z^O_�a8��?��s{}��W}1:X��q�T�#KpX��pb�/CDP�f�nݜ�#�qq�8��۲�p�!�:���} [�:S��.�����y�2Hz���3]�#P���K'�s�9[�?���s����n�����Gu^z�E_�������9�l��bϽv��휰�h�\���.��R;��?��;��KN���3�x�M��뮵���7Rv��9PJ��R&v�-��Jns�/,��_~+N�f{���Χ_�g�ζ��~�+4����M�3����l�~a%a2���(T�Ē�p� Q��;�"���:"�9`���=]x��ܬt���d�;c����i�jol�2~b�-�EK������>74�Ƞ����92.TT��2����(�(Z!l+y+f��9AL���	���&��(:*Mt�0�Ǩ{�X��~	�_P'6P���_Gp�főN��|�	|@S ��P���M�m�Mf�����('�Ͳ�_~dm��,?Wa��Կv)G���묣����>�l������c�k��f�刌ńY��w߽�\{��>2�-�!��n�ʀ��6���fn�������#�Ȳꚥ6SF��ɓl�)����%�%ǆO�٢����6�|�M�6Ͷ�z;�{ۨ�V���ą猙3��+.��^}�5k=�>�&��A��7(\2�p�#
�(`���_\G��0�9~��ab��4����㼃K���4b�(�b:@����џ��!<�����?�8@�g,���}k��
����2�2���G���?@������V�E^B!�����L�KH)�݈Ϩ-�d������Ib��%�(�%nx睍�\�J\��6�Зq����WO�-c��,a�1�,_i0b�O�����aC}�{z��c��mԈa�L<��s6g�l_5u�T[*�QΈpF�y�?�w��;F|j��R���7_M�'�xR�ʶ���if�Vfn�������I6j��t����Εl��&�HG^�5VP𝥊3g��%S�af����x��"��}��o�u�jBp���h��/��'�zZ<��z��nS���XړAJڋ�߼ɗ�R�B�1Z�`3
��]wݥ�&�"{��G\�ӆ�}��S3��x�5���o�Y�4��^{�m���i��}�>�����v��t�)����<�G߾>[���WxδY��W_}�4�s`� ��/�Bz�2����;��2\���˯�����ܠ�SϘF2�ޗ�h=b`�><�dfg�M6�6�������Y�����ox���#]���K��ǉ}k8�*q�믽�G����[6f�wcΑ������Y29~�W~�رc������O����u��������V���2����~���_���������j۾�=f��sf�/).��	� ��O���'�9u��}5�2��jC�q��Fp\X��x<��K��C����C۰}�2 �ӌ|"�!�$>�w��p�3����S�ֈ��T_~@���W�^ϕ�����9Fe�z����Rqq�J��w�>YE���̚�E�辤/e �>��D��%z�K殿��O����0)�D���^��E.H�Pç�(�� ڻ�_�_kkK��1S�.Bl��]�q4ɿM�S__�����,�(em���{�bF�@@(	�$�lYk�2[R\���K� �������v ���8#R�!>V9�0N
���F��%2��}������{\o��z�b�r�����4[e�]��
�~򉏬�7w&m���/fS�N���wƼ%��y�Q�SyN=�L���K�N�k���#}.��"J�Bf ��3g�ɧ��Ƽ��z㕶�����<m���em��b埖�+CF͐�QV�٘˲_��V� /���z��u�O8��G��o����H�)�#|s󲍋E*���̳w^{��0D�\SM��
�����Bk3>`�����a4��+%I�-�?ύ����@/�;�ʨjaQ���\�����c�ͭV�p��4���h]�iQ��A>W�+��􇀥.�(gT�g�mjV�ZD���s߀؟�O}�(�E�0� G'�P�ĵ�o�OkU��uV��n��-���޴go�ܚ�[Qi7�,���j�B;�#��n�e�������B�?'*�σe����
�b���R�%)��`K��)���#��è>�
QII����!`B}E���~o���j�5��ؓR��Γ��H�L�~ǌ+Ke�8������3�<�Jٖ[n᧒qd3e�isA#˛r9�����3�IV(���\@�����} ��NW�H#�2�X�>�&��О<�0�[h����}A[��F�q�@{�It�o����c�W��X�����b:<�w�1h�E�����O���u��P�d �V���m�}@"���쏰��>Ɔ�{�k�d�w�]�{�PN��%�K-��@�ǥ](u�a�6�gס�A��*.� �eW@=e�NK��e2�j����ZU�qg��Y��o��3�<�>���0����&���E~��p��%G��K	~�E��x�}���A��3�w�2�g�m7�6��ԭ�����:ʕ(x����Q.Q�������[o����)���Yz����Zk��ᾝ0�~��N2g�������X}����=w>fGu���m����Ϸ�~{?.� 9��d�a��� �jkj��w?�\��싚2u��kw�y����=�ǟ��}��ߦO��v�u��fS>��4��/�J��m3�Ou:���{m��S:�;���;��Yn�� ����J*�	F
e�o�����n֫W_�l�E~(�C�|��}�}��f�����h��4{�*e���^v͵�X�L�p���n��OQEv�N��L�������_(Ϭ^�^t�Ev��G[�R�f�W;��{�[k�$��E��z�L�>��x�M�CX�ž0���[��ԋ2�i���9�e2���!/���t/�e[Đ�C����t��u��{U���'���������X0q��7ݾ�o�~��.�mUU��%�u�/x37M�y�Ȼ(.�	e5�+m�(��#�"o�=��Hc��?�ż d�B�d��Ѧ��N�9�oVN��9�E�X��Wh�4I_<��L����N�m�_� m--��_���znN� -+����^�ꫯ�������o��_u��&J�z!k�0�����u���c;��c�c
t�]455��"�B@�
���󟷊*��.a��L�#_�'���xii�J�1�����Ӓ-�"M�O���Ǽ��#^���,�t!+[�S���j�H��ъڪ�����G�yZ�·766�777��]}3��]����|��J�ˤ̉�Pv=��� ��Pmj�+m#G����ʫ�U�)7.cI�]OQG\���O?���[*M�\Z���Q�Ath=?@,t���г��²�C����8[m�U���ǆ�d����\�e�]�P�)r@/�5�QY��y��}ח�pQ�c�?n[o��r	�8��K.���7'�G{̶�l����l^�7��I'ەW]A�?��]v�epk�)��n���r�w�~m7]�m��Z���{��O�a�<����J�HWK�p�5FG�/'[qrQvf�1u�f���Bɧ�H�?L�$6��	'R��#[i'n�D9�op�����c^x�Μk%2l`^�J�b� +����K�̖'�����w8�Y�T�&O�TIaB�`��vf��ўP-�쫏>�態-�Y
�h(�[���ݖ�߻ܦ��i�#�����:h��!�p,DsBVW��q��$71F�wXj�K2�����˞#_�(����Tk9rg�nc+��k'�M���u�P{*Lsc�U���~��t#RPR���;唓��;�r��X�t��0E�H>�.��'��!V[mu�)b$Z�O�,�O�>��FQ�5�aƌiv���Ҕ)E��_��?A�ׯ�[o��/�ʎ8�0����~���+%ď�ӷ�a���������b�"���z�M�0Q8�@R?m�^��e$N�����8�юс��'p�#���0|���>9n���%|���;a�b���0j�/i��Ox�4��	Ź�q��8|'�2�V,���p|'_�S^�c�q�z��%�����a`�꠴�����e��ٸ�]	���l��ֱ>���z�)�l�����X��2O���2�Ox%5P�~��S1ؕ��|�S<A��B��j������s�gC9��S�8e,[|�FP�(Kl;:���:�'ڊ��-.�͖A��2��2�R��U"#����h��l�mm����ϳ�mF{%�N���W]k7�p��ow��J��=.9 .��q�_�@���k�{�@zT����7^w���m��r+,�����s����c���p]#B�,^T)��v�뮻��&�y��W�]��G�Ҍ�3�@BRP�c?��� �?���gN7���WҨ#}H'��~�m>C	Mq}K4�h��s�'��׮v��G��o#F�d+�������*��~�ls[����F�@l{.\`{ﳧ]{�VQ^�er��T��$h�6�E�zک����Q�窿f�7ϱ�;�^y�+������V[{�u�D=�{�'L�ڍ˵�Y���UO�w�ʌ��0��[oټ��m���aH���_�6a�6{}{J-Y��6�x7�	���nW\~�t�K?����:YR؛�sf�O����������W��%E��K�Dύj���f�OԐ���ƜtU:��'�##mɒ%i�i!-]�!~ฝ�m�3&��0S�r�v$>�����վ�}��אy��D��FW��<�K�%3y�Q`L�M��Ҫom��-ʫEi�fee���~�7WVV��z���ҋ��׷�G�&S��ʺ���������ɓ7x��Kz��QP\\���о�-W|��G���W=�г��LL$�,��ϟ?�P�&K�p�̙EJ<OH�@�K �e�R!b�d+����w��1���3�������BR��אqy��˯º��p\��%?�[�"z����Pr�K��h�euJ�vqV���6�pLGe@�';�Ҕ?���H��-M�bi��S�<!���l&�ԣ�.>z�_�x��i�ccyyyu�>}Z$�J����I��(��{�N�:M�g�uﮎ��c(ٌ��P��54K�k�W:A� ��L��o��wr2�)o��hBΘ�Q~L�s�rmu�yo��p�����"�M^o��m@߁
��2��}�=`��r�w��N�����W_ݗ<P'f���v[W��jʴ����^����v�Վ��s�r���yv��g�ŗ�v��+�������|��f�w�����*k[��^����������_L�~����^R4�����tR>��ȑ��������E-h���04y��!����>E�߄�bF[���v���j3�@Β�[�+!5w�M|�mk���]��Z�|���
	��K�����Q����I�(PY�ԡ<�)'�]���7f���s�g����	��GF�+���`�4�K�?�;K[RcV+�R�ࠍ׵�k����Fu4�]�C�1l[���J(%^����紉Q�|��:�@�H�s)4a$�I=��]̽�ں��,���<m/�q�H��rD_Y�R�lɂy~��u�\�o�I_u��v��O�n%�n ��(�(��w�|*˒�ň~�V�n��=�˭XF&ˊ�{���#�,i8`���JY���i2��g�y��=��n�}FW]}���Og��7�����hg�y�}��D;���|��#�i���*	��{�ˮ�v���7Ǩ��,[��RP�=h+S�/��),�Q}���z&;�*��_z���3.����p�H΋� ��w�cY�!ƍ�q���;���@Z8�BI����cSk8!,�|�ԋ����w4��0@,J{
Qه������o����\su�ǬW����/����_t�]�m�Y�fKAQWZ�s�Rl�%N\�=Jz��rJg�/�n/������c�l��q��)�
�#�7��b�QHkj���w�s�����rC��G��� �7�&���
�Ώ���u� �_ҙ2y��#]F�C��>gt�����a�J�lM[u���N{��a��`<��j���
0�o��.IW��5k��~��#��j����v��fϙ��V�ӧ��G������;���>V�h��i�*�f�M6�D}���ee$d��k�� V��OI>�'e{���R�r�;o�0���p�����Ysl�С��b$1E�#M��9���;Wufi�Q�/�=�����1ʝX%�'x@cS�ډ����m��]v����ﬨ���[C�;����_��7���n5�5��OyX:}Qh�>E�0���v���~G�*eZZU+9����V��$�|��:�����.����~����lGq�����zS�Qt��Yohau[�a��<I�-w�q�
��Y"�(����x��ɠL�Pߗ�������9�`���+� �9;��Zw��vO^rɥ���]��}������W^�G����?G}�k)�3Է�jk�$'�ϝ?����\�Y��+���*��!u�)���^zu{z�~}��R'zi���=e��l�i�j`ώt�,��L���Ou�0�4H�굋�1@#	M��EOY�!s���d�+/��A�f�E�1�R�y�L5�	��5I�։&ke0I%lhV���S���U�|�f̜���܃:��#?p�#�'�sϿ�}ڴ��Ϝ6〗^zqM��Dye	M*K�\�h�E�+���ra߾}=���p�����Ѯ~睷�������;T��xg��d*� ���-U���\$F,)(��[��)�4:/�P�m �4��i�!ɇ_%�"m���;i��w����ap�ya��K���@�)).a F/UN�d�`lj�7�aԍ}3LU��c�0�����`aCk�!��Tq�;'7�gU8m�\.8G�7�kY��,��0�\gH\؆PB����`��Qs7/��M�Y��z]���t��2"��H}��
�,�IWV�R�%��Iaey'�[i���^*N�d<h�RH��~�N9�T�=s�_w�5������꫾	zx衇l�m�q��r�+�*>��8��G������]|���G�r2L�iӧ���?gw�q�����������5-��es��ޯ����l���W��hU�;x���xiR[�K��U�s�{a��2V`�-2��}	<���/]^5�xH0t�[oz��55�~�5�!����D��5.�����Y�܅j�F�*-����be�{�l&�T�ڂ��9�[1a�p�	�R`i��Jqn.�3G�*ߏ�fʎ�N_Y�#�-;/�*gα��b�S� ����˲k��^k�P��6�8_B���c�!t�*����[�.w��K)�Ĳ6�3�Ğ+�j���9m���OI��Df����ʆ�Za�{���q�'�=���Y᫾ƪ+��'�hW^.�IiW_s�����-����=�o���[ǋ�o��k)n�)��ҟ�,7��1���@��>J��D���
�Ψ�R?*�M��ՏQ��4߫W�A,�c�QH��j�P����<o�_·�^Bf�ω�\ʬԛ��nEE%�+�YsNY�v�"ڛ.(;y��Aԓg�?�_���?�&O��v��E�_�#߂b��&���g�L��&!]ʊ�i��:0p�1�� y�4��@����G��e O\,'	<G? ֑�<��K.+.9��DC(�l@A�Hao��[o!z�����ܳ���đGa�gL�eW=˽�$��p��\?�A%�=zz>?{�����| �q_�b�!m���1��XL�Si"0�X:4o�\�ԍ��&N�f/����z������Rg�������dP&D��p����|��Ͳ�ض�|k�����AR{�.��%>r����m�-F��ma�+�������t�)a	�m���F�W��%v�@����l��wu<�����c�>&*a ��⻒O��R��"��d3��\J
��9�pQ� �)`��_���7�|��`�H���n���ٿ���G>�D�sz3<�2��Ñ�#�F�<3�3o�l[K53HH@��������[�(١���P�V�9��K���j�3{����~(�ꫭ�rW�&�n�/�o��@zHg�x'�8�P ��rlv��,n�{e�UMҍv��v��׹~@�$�ؑ:t���%�:@t@]���_,�g�=�P�׊n�x�����M7ݢ�����y���fN�m�~������}�E�|��dy+������:�n��{��?ޟ�����y%݊l����c�=�uC`�v���k9rгW\q����e����؏��y���{l��Ƌ{��Pun���h��oʒ.�WY�4W��`檴��E��&��!��1cS�Д�p�B��Y텅Em��[���t�!�S�����v�����%� ���C�TO�����Pi�-���A��z=w^�0.ٿ�v��8�[۳�3�JK�,OTsKK�t�֜�l���V�q���ΝӖ�_P��>����]�W_}����9s��J���E{�~�fKϕ�	7�N�41s��yM����]v�ea"������ٳ����C�8�...�D/b2�,˸T��|JA�!p�;�3���� F�������.��8�����#.�3ߣ��72qҍ����w~y�<ġ��?��_ 8�ɐot��Vxa���*ld%u������7��3���rI�0K���'AV���c@�#��%n\ �MϤ�;x�E��<
]����8c�~q0|F������GE\����L�*�V`���q�,	9���d�n��6�,'�p��z�-�HL��믷�8��_y�57��#�T4�ȃq�Č|�A?����������¿۞{�c�^{����p���ҡ/��b;�lf���ۺ�����垛EVX��>���.��q�Ln�F�f��Jk�q��������M��Fe��P��6��d�u�;�tzDi�]yD<�M���/��Y�`��M�J	�^�X��	
�u�^3�e��wh��V ����2�
�̛km��YP�c���L)fM2*`P���X�F�0�se<L��0������j�2�
����2n��.��ޢ:�ڞ��\}�����tkHk��=F=O�B?-���$�2@��Nj/�y�:�4�i0�jk��RY�=ӫ�{��E��a�2��1���`�͵N:ɏdŐ.��r;��m  ��IDAT���d��[Yw.qK���,��c���R�'���ü��J�d9e",�} ��Ϭs���"�b��K\Nsd cа�����Ox	�c8af��'}��w����7Ǹ �gy���̴�8�W���q�^v�H���!��p ���W�a�G���B�w��;
H��?B�&�_�>�$-�	����G�&l,�w����1>.~�e��=��b�����3�4���4(7i�A.�H����{,+}�e�{�kܭ����`���^�ܒu�
f_ã�=�{I�/��
���&�gCO��X�����)��1�An�n�ώ��`~Ю�K	���f��*t�r�����\=;0t��%��B!� /�Il��G��0��	��f��=l��@���C���uv�G؎;�j�F0��@�#	"A&W?���G�;�N*ݠ1b�|��*�{�q�}�3��fL_k���_�x�~80��Ÿ�m�=~c�gN�^�z���e�}eD���~����s�'��s~��1��f/�����ܘ8h��6�=b�/ϴ	����!6�5t� S%=�Y���%�͐��Q��4�S��e�q:�7o��ǯ�D7�::���1���ؓO<%��ź��ZV�dA��Kt׷� ��ɗQ�r�/79���-�;�8��'�Q]�`g�y��|�M����ƺ$�/B��v � �.]����o���[�H��ꆾ�.yPR�͇-]�KX^!���dU�����ś$���;}�~����,X0OidYq�r�F�,�%<w,�.}�%��J�ݧ/�>�1}�d������?饗�RV�c�X��A�kFKkKZiIi�"|��$@/K������>=z�(��I�������q��B� ��A���	O�F�g����4�F��##,P������2��o<�4H��(�����K�NfϞ�kN��"oʁ�\���K0��?a��m/%iᢅ^�X~����ӄ�ρ�0ȗp�Ɉy��'���c=�eG9�iw|�h��: � ���� s峝��w��C�B m�aH��&\)Q��)_��ŗ_J0��M�[l�����V9�x���}��_�>�7s̱v'��R@��]�eT�uFT)3q�/Bߕ}���`�:cVڔ����N5�!�%� �@ ��{�-��B.��1+��o� [eݵm��+9C�c��}���b�`�3�Eq�Őy&��RA�Xc�\�쑗��ɐ��U�[��a6r��l����5��؊z��E��)�a�r���T,ї�˻�_��p|(�0z�,ĺ'ǧf��e�_m}�oB���{X�t�i �
��e2@ �B�
o"�8�� -���E�L��9�I�c�22�0d@�c��O��q��-�l��e�%R�m�I�-�V��M�,����7�B��fI��8m��NJ4
� �8�]��p �Ñ��=9��F��73��8 �.ԕ~nȇo��3�����u��u���p��|���/�,��<SnҊ���HN�?��C�w 5@ʿ�!n,;����D�y��}���e���	U�U��k�������3p�X|ލ�|%ONBd�2�"��Xee�f E�8�%�L�3����Ɏ�������ћ�/3!�G���C�x��� w(|�K���?���T�m"^��8�?4.�m�}B�^�w�C���_|i���p3���I�T!�n�o'���}y�1{㵗쑇.��=.���)sP��w�݀�/��A�rJ�����2���2�d��^"܆
�A�7��d��/������ɺ�[��z���o���)��)���?�b2�w�E�_|�p@��b.gЅ�V���;��z��r�@C��K���>����s���lx��o����'�Q���z5C�,\�p����e���ˊ���=��.���e��n�{���(w~O�3�S���.��A�F�AO��#Gٰ!��4��r��2����)c��������F3ye�9䧇���o��XI �g����@qJl��6|� [c��l�5W�!����!��y�UF�u&,���vX��Y?���L�&Q~^�W����֟k��L�g��+&���zGtv�*D
�GY�! ���9��ßw��t����a�C���<�%:!����y��� ��o1m��Q'��8:��Z�N�(�Y�Eq�L6�Ó��Q�Èf~^�!�N�r̲�b)�"wCa�G���G�% "�`��K�)Y�EZ-��.��w��@d)�Ǖ��`=���w00bD|�@R�Ȱq�]q�W408a��B뭷�3��_��"���r#5���.;츣����� ?��êK���O����}gw�y�3��F��4(c��M.��`�o��������z��.�o����]w���_��PZkhn��Պ7KJ@����51���C�1ᾍu�bYG-�6*����Gn�/����8Ӈ���b�r�|1�P��#^�ִ�_2�ƌ�z�	��D���[�e��xG��Qid)��2�M���xl����(�^���t	��<c�-V�Pg5�{���++	9\��Ҡ<�)S�v�צ�=,uT9�ЅD��/ay�3qЁ/9ٓ�Weʊ�Ֆ+[VC������*��헽�pk���ޢ�ۮ?cƼm�����#�ٟ�2��Ж�!m�݀T}�=y;�K!`�NuU��!�Z�]c��x��g���TZ<�ɕ<f�0�����?��/�|��)~Td0��CGx.�$ܒŕ�����	�n f���xh� �8����!~�#���M�}!�c9��я%�����M�X.� �c��@�O7��1\�qI'����ȓt	!��_'�S� ��#�x��-�=�ۘ/!o���������1D�{6�O�r�ah�8�p\�A�����A(f�Q�X�	�f ����%NLYRPP(>[�Y��@��R�.zE�E�E��3��� F�����'C�I�38In;�23�l����B����gR���zp�-�X3�N����^x�y�����q���}h�>�=��6}���N��أ�>l�\r����{�)���G�w�y�jj���iѢ�3p߳g8�g�̹��C�� �j�7t"��3�9c�=���V�P)ó�p��F�G*m���.˺���:7�8�y��K/��O?��?��3/F�+�����/�qVb�+$0p��Ӧ�~)�2D�E:�t�!�_�sȌ�TY��k|�ۻ����VZR,CA�ԽL�)�A��s��ho��?��C?��:`$Q�)S&+L�t� �k����`�U�(w��kz)O�u����%<si�/��t?���c]��T_� ?��,MeIj���������%�T������ NDX*Cy�	~�g�pY9���g%�e��XZ�^�~ ����*&L��u���d��6z墋.G��_<tJ��A'LԈ�Y���:���v0���B��'N�pf����p��@��.:u�E\�|b0�q(1o��!=$qȓ2GG�0�֭#4P�g�=�ň.更�)
#~1�PL�VW1ӵ���[ ��D�Y&6BJA��T]�B�(��z��Z�F�XVפgF=`R�Kyp0Q�12���)lg��C�����_FU��q�1�[D�M�%\����mȷT&�+���3R�:w�0k��9�OVn�u׵s�=�N:�d;���; @�(�]T�'$l0�؇ő���;��:J�.g��:�{���8Z������v�i�;B���I�V���UaE��ߥ��^f��i��#�\]�w�H/���nY���,��L�"]����S$#�Z�����'����Ȕ��T����9]�r~p��R<�K�t����l
��LP���a*JKu�#�G���V��s}I]#{qX�p��F����#���oa"K���8)�ц�)(���9���{٤iU����f1���V�`��"v����~��0}4DG��qO��K���Y�	]�_n���_�m�Î~d.�3ȟ�F��ӈ6���@�Sd��3��3#�(��7�U��$l�gP�~Υǃ�뮿�7C��w�9�\�����S����'�Ї�'���I�|v2�(>��o��?���s~��?@ZQ&�O���b��<5�Gg=I��ģi3~C{��8�c���<G��e�q��b�t��?˄?�q�<��&Ə��]o�1˲�����C.�j"���b'�ygT�,�[�e t��%3�|��-4~��R����8XyC��;���s��M���S!❊���\��z�����?r�%ӫq�X�2b��;os�����`z�n��f;��c���%�,�f�7{���ű���c�R�P��I�}��9�L� 8@nbp!gu5{��T���SN�C=̎=�x;���d0�q\����������_��:�����>���lG��"nG	�/�9��=�=�����:��q��/m��S�����!hnf@�%��2b*Un`uO�͞3���a���Et
���Ch�f�d2�6�@�UZ�:\��;�ĞfX�"Pwp��Q��e�����o'N�Y�g{�+�V����|���3m欙���o�	�m��q6�ӏl����)g�~'��
�6Ћ���>�1}��-g�����%l���6Cqgϛe�ep��I'�!�^��:�#:�PVVn#G���}{7J�Y$�N�\�x�A2�7on������d���D R����������t�(�xFi��3��2Bg&̘8�!̌���aQ�;�"T���X̀39��/��TvN��HD?^��H���9�Mis�^{A~~z���.���Ҭpl ��kmQ�-R�y�,�YY�m��y~t��{��l� �3'v���Lk�����l�S��3�đu�����zς�"��g�~Q�;e�~g����P�8����&	JE�8��&���oܸq�Gx��]�Iv��U�d�M��V^�n���`�u�]1O���[o�6���s�Y��C	%�C��{o7d�~�9|�����Kv�o��^y�Uv�o~�%D�8�3�+.��O<ɮ��*��T��c�=�#[�,��.>�|����ګl���]~��M\�d�����<~��f-9%R�E��W�娪�4f��y�g�p��� �d�K`�@�A�qJ#��2AQБ&���I8oǒI �����#�IP*=Q�̸t��ͷ6�s�����r��U�.s
r�>��=�̅HkIdE�^j�I�h+TC���Xn��#���6�K�oɶ*?_ާ�22ٯ��f9�IE	8���E�1���8��}Z��	��ʃ�q�w����i㬴 K8j��ѴF��l��	v�W�+����_h���G�
7p��a`���{ڌ����6%i�5��m���}���A&W���9��#=#�ψF?��C��Ȳ��D�ry_vv�/ǡM��e��:�7�/(q�c��H����u�]v�=���.��ۑ����`"�g�z��2s�-�7(wh��풢b��g�u�q�-oOe(��x"?��e� :��/fР�H�8�yP_ ~��D�F������Q���x��a��f��7�ő.a �c�@L�tb|�wh�^tƍU��"�S�2۽�ۋ���ٛ�>��v�c��H\���/qI�|�'ߐm��XF���+	'���QD_C΢�1�F�7��r�!^�/��gDTj��#~�]���3���㦝x��'Cأ�I3�8�w�۴�S��$Ǟx�q�t�p���7�c�{�轛�O��"Kkj�n��>��3�*�1�Q��K�7���}����/%�][��B�S��RO8���p�M<�O�~i{챧�fN�mS_?\��*sX���k��o8��͟a}z���P3N�d6�<0(���A����7h����2�CN#��(���>���x���o��a��0��o��Kn��FU.��q����ng�\s��U�/�!.����0p{�5�����+6(7�3����:�^Q��㥗\j��O��x��>A[��WY\w��v���y�:M�z �� R�tB�/q9�#��9�}#�#,�ej��&fQ��H�S��t8}� ��g�"�i|	�c���!9��<(.��1-$Nf�����۠�~>�v�}��ǖs����on/)鎡��`Y
L�/���b�G���Q��oh��MrU2�je qP����BH�H!r��{��C���D���(
�,ب8�A]Ȫ/x'�0��a�L�#g�s����g��c{�� ��`�XB��nW�k�j��_u�j嗱dɒ1�B��UzFz[KSK���K���\�XQQ1G�]������ઔ+�`朸ל��զ:։��F5$@��	�
	�.Aج4�<��BT'̔��]J���=U��o)�k"d�us��+�Q,F��[�Ɛ�r����#�P�|t%7�@�9ϧ��$�9�>ю�1��>}�4�|�{�ű܎�y`�e���&�T��oi �G����A���n��Yⴇ����O	fS�;������C��#}��,����#̛9�N9�4{���즛��mw�٦W+�^�g>�k��V���|`�?=K.lFu+I�1���6ǽ\���`Y	c�_x��(��������yS'�rǟ�)ɸ�@X������>��]A-,c���--�h�"k���d��s�Ag�p)���y֐8��n�(]������@u�pИ��W���'I�"���l	���''E�$)<p��~-����;�A=E��8������� �I g���琉~=l�W�ۧ��a��'XNK�p�H!#�5�x�;��C|�[���?��z��F�}�&H�\�(�2�3������ͪ�+m���v�g�($7�c�pz���+f6��F���U���X���+��U�!p���>���ѿ8	e�2֩.(V��>���	��ex��e ��郜V�w�!���+�$�w쫑�"���H�N����?���t�闣��)<�x �b;����� ���y���I����CJ�|�qx�
Ϸ����p�.������x����0��3㶤r�͚9˶�vk�GR��}��^���>� _��+������.���W_9?E��^8,�Y#f	0�������Z��?����3l���n�1s����w`�6�N9��աÇ��E�m���@t���2��U{U,�1:p�(�0���A˸ɓ&[iY�=��#���@�뮇�#�V�2��K�R>�Y2P��GZ�5i��ԣ��Q<J�mV�J��ѧ=�I�Č�0 �%����,���{l뭷���c�k�}l����~��r�-7)�g��v�	��o&p:Y��@9����Wů�X�4f[Q�H�:����X���-����_}�M�o���Sk�Aħ��}����Lz1̀�p�4��V[m5[i�ݐ#>���խ8�W�0���$�U<���1�1�1�b����O[B��*ڜ��&���o9~��СC��pJ�_�,����L�:��I?ʼ�h��������[�u��78��A�F~� IPGR<C։��AB�jZ? ���q�9|a���X|��G�e��������PW�� ,K�)���N�>��:�()�k�SP'�P�߿��Ç�&&� �6�X �t9��_�O�8��E��5)N�:��-����0��8�{q�F��e��{�r��:�w�#��x�\�J�Iy�>�PZ�@� �4�NxAFsSs���ʼ%��R�����s��*%4�S�Y6��@Wac��
B=q��[J�]4{֬,k�����b`0)!�Aeu&�H��9�:}�͝7߅L\j��8>a�(lUK뭭�ݧ�:0�� F3�`rÆ�!��5j�O����3;��ꫯvaψ�z��K)c:�������w�b���~���o�PN�a6!�T��;��R,���������{_;��m�������z)�%�~�!{��'�߀>v�ݷئ�mgc�,�s��׾k*�^#ױ��k�<m5K�0V8ПT3˔ ��Z��H��^> �RN�%;	�*�^�;T@�!?f��s��z��s�Tm�U�_bi��2�̘n9%y��Zk��3l��J7vhW��@j���`�\�	U�}O��*�+}���)%�4�Apz���i���c�qi)�H�E�,S� \P~f���	$��|�cp�;���BY*k��u���8��l�o\d3�<ms�y�Z�α�\���Ɩ,�����������_`���e$�F��%8���p��'��C���!��N;�ʗ�2��b����L�r�UV^׆�)���;�B���[T)��,����*z���Ӂ��i�&{=��d��hl��V)"`.K�
NX.ʑ����_|���0xY�	� �F�ڔS��r}�����Hk]�p�mp�ߓi�~�#<��N�K}�i��G�׎4c8���@��,(� <���sޓ�� �ĺ���|�?�W�I���2'y%�`ƃ�أ�B��hwĭ�-�����.:���ݰ�!c���>��t�y����`��1
)�q8y^r�%6z�h���k�dB/�ZY�ϙ=Wi���ٳ��/��}�G���.R����ǟ�)f���@I����q��c�>%_�'mK�����%�9>����a0��^�3�8K��/Wϊr++.�|�m��VB� �v��:�7��1P��a`` ��}��K}��;��&}7�~���������w����B��f.�?��,��~8��9JY藼G\7���6p��a��?b�8Ä(3a��O�P�ǌ__s�ʳ����h ܒf�=iy�$@^\}����~ W�[�b�v��bذ��ߪ�jħ*���u^H>�ԍ��~ÌMZF���G��,�oPݲ�����(X�r�'22�����U��K��(��[�Kj�"v�]���@��`�~�-��n�c运��� �'�w�8n�;A�Jm> _Z�qџ� �=�]l*��H�oa��{���+d$]۽{�JOd��!�⺄%KeJY�6o�<f;�JJJ���k��y��ou̴���#����s���h�TKaCut��L�����#�l�e�07Σ�U��9�m�R'��Q�����;�م��i3�ĬFyy� �{1���;6q��v�}���O:ɍ9�Ex�P0�"� ?�X�4.^�H5�O+#Ͼ�����Q�L�D]a�P+))��0��.|���z��47Y��$�k����5�����;���,s��6t��mqS�∹���e�4���r'��K` <�h��D�R;��p��RHx% Fg_� �ַ&��"e��uHl(历\FOk�j�B�nT��f�=c���*�57\���R�X��r�����x��0ӣ���5);[H�_�UO.e��V��s�8P8�N�fm����0�@y7+Mڛo����0�Z2���A
��szx��|�_d��3���O=h�i5�W��L�����������W�.�V��߾��%�%�`qr��=d�o%%s/G�3��q��UiY�3Ψ=�GIa?>l��j�^|�^{�e1����؈�C���آ�6���RTx(TӦNsZ/���EJc�M}f��G�I
Ǖ�Gs����o�mWm<-�?�y�B�(������`	���J�"4�[Zés�qS�p@L�#�D<�IG����� ��=9x",~1N�c,O�!��_��-q��b:��
�?�@��g��������tֻw/��_ϳ��Z۞z�i;���}Ч3Y���!>y����Ԭ�>���D�1��b����9����Y�X�4��BW�QZ�|��������ߨ� �v��]m���J��n��?����ã��?죣lG��ଓ^H�>̑��_��z?io��x�لof�Y��z�M{���e��DlY/�����p�8�,�/������@�́��f����[��s�**z�!�h�{����̦�����AnO<��J�j;찭=��?eȔ��5�WȀ�ϩ��fVߏ��{p�}a�$iQ��<Qw��� ��	�tK�`�9��g�}�.�}d����x�H��4��߀�i-^���
��d3�p	.4WV�]�"�\�X�Yo�`��g�����˓�������Dӹ����#�KK��~�����(�=g�-���������oZX*�s�zA~7�7�d�(?�ܱN _�������@.��IZ�?���>i73R&7������^�X�	�D�N�U��?�L\�.��}��'�p��'�|����]^J�~y�B+�R��]t�E�?����*-)Ƀa��!�83Htq:)���Kk\YD8��*�	#�@v�J0��������(y`�ۏ�V�g�5b�S&O�1�c7�x�����HO��9AI�;Q>'_e:�`t�#m�)�7#�U�J���|�'~0q�dS�B�c�
C�y���B4��1I�y2��o�>�����F�����i\o�
ذu�����b�RZd(5KC���B��x�b�,���>��h	���e�[�J�e$�	� �u�����WY���0�?M�ono�&�헱f�[C[��Rlu�նd�\ˬm���6	�Y�?���X}1f�F���#[���(�ص��o���*$��¦e�,)F�	H� �.��]eՁ�P~pA���;���ѳvڂր��"�4U���e����3���n���<i��$���+zh���f�n{�aw�uW��t���n����{��a�T��7y1������a͒�m���?�0W*9�j�fjY��{�`���q_~�57rpB��@�hp�M�������ww5j�_~>�7t�/��˞8�h�UVu�������02ͽ6(0���y��L�Au߽���Z�:�R>��+E��,o�g	m���Y��5pc��B��p8/���"�]y�KYQ���	�1�>����[lcҌ���p�7}�e�9q�B?�Qx]��O�ԯ��*~�E?����(���Ɩ���P�X.�%�ĻCHN?z m��9GmEz|���ť��3�m���ٯ����t�v�(hF��m����[oڻﾣ~��6�t)���w~�;�y�m_��λ(�&4�[e�>��}!Z�ۧ���6�7���c�	�ۏf^�De,�ztʅ���G�m�A@�~�+GG����g�<��������c�?j�n�#U&�L�-���'�xڸ���>�q�*��K)O����K��M�dM7���`yآ�%�j��RJң�����Z������k��ћXqq���4��/�ĵY����6��2<������	>��y���M-n,��ya�o�O >;�i���8�M��h�ߥ����7�\2�ȗr��5�\k�����aw�n�m��]w��*zuw�r�Ƌ/�`K+���&ː�+��e�o��>#:b�Jֽ��=�P�j��9ַ_�t�A�������T����/��M7�j����KQ�BkhfEJ��h�3'��-�/����]��������)H	��]�3��p�U��'�!������`u}���
��-�?���SN��SO������D�+���+��_pA�T��k�mٽ��ې!C�#�ql(���6$r'K�����֖.Y*E.��W/��̌,�Lϲ��Z]M�+O��� �;2_�c�X��쌚c�0�4x�@�D�cs)qY��l��ћ�Rο}������H��-��I��Y��Z�����c$�io�8�0 ³)���	#�n r�����É٥�Bf�
�����*��K��>�J��m=�ˬZJÄ�U�QXj���V��2�U<�.cS��,���4)����QC}MW�,,��A#�yDg�pY�/�bd>]i�e�Y�=�v��I�-T��*�WN�mY�M��*@��;Kqkd\.����2յ�O_�Ӧ�R�3������H�/�%������C�HV��)�(��:��vF��g�T��0��_���?�x&�/9 9՝�fG*�R�RB�(I�#S�a�o��Ko�h��bш���R��.�A��e�5��%˖�kl�UV��v��G���Ï����(.o��97V娲���+\pb��~(P�'���K/�,��r�t��[���h{���ts�n�?v�5���-��ʪj�W��zyV���,�4�;[�h�M�4�������go�5VM���k����_y��sɠ跴�m�ɦv�a��l�����QcA�vb �G������]]�J��%J�6U 8�*a1"��_�{��'Q����"��#�#�V���2y$�B�D���K�|顊� G����̬b�@S|���1��Ԓ=s^&���3��/q}�����< � $�O$���v_��_�wN�¨��\v6�p�|_�i���N��^{�)et[��9j��`��N2T��2.���~��;Ȉ.�w#�4?��2����dL���{>X����^{�>��+�!U,��$|2��@ �2|�U (۬,�x(�,�Hb�ug�>ԁ)���9������s�-�4�l5˯@eE�
+��X(��xy�7��1�v�ն~�3��6�c\���\�`�UU.�,����J�3o���S�t��!l�UW�����?�p;�ēd8�d#G�����B�N�<��>����ۯ��aCܘ�6m���l����(9�A��F"u^�7�,3K��!Ja�Ja�r.�*���p'��%Zz�A�q4�O>e�s���{VT(��C��(��H�]W�������ϝ#��a_|����:��WFw/9b��L�3g�+�'��x;��ăַ����+��dhn�٦֣g�}9��5k���^��pw��7X߆(l�^��j��.2e��v���O:S���=J���D�T�e�hw��Jo�ef�r����_�W���:��\J?p��wIy�t$�,Mr_��	�!���M�a������E��4xf`�l��в/U=����X}�o6�xӷ.���p��
��M�~A��ږv�=�nw�Yg]'�8��)�l���¤(��2ȕG�V0B�>
/K�PӤ�b���X��d)@�s�<� �Yi����ڔ)��ɱ��u�3�M��.���$�-���
�%�*7T'�#<`�<G����7\�K�0��0����t�I�"B��T�Gn=x��ӵ��hw?1Ʈ|�#��?�2{�EK�De�P�$Ó��j�q"�?µ�cPep2�������gJ�Kf�ޡ$a�<c ��Qi禉�����	��x<�te�+���]R�&|k�Sf���J�_�V��4��I�./�a��zF?�	♽[(�1bF˗���� e��?j�
K��`O�♭�Ap	_�,��-�p��j�@jK}����:�ݫ�J���;o��_�A�--[J]M���U������ �_y��v��V\Z����c'���\4��q8Æn����9q����~w��$l�����>Y�}lQ��K5�9/T\*#k}��[b�K�Ϩ/֥)��R:{�h��#��зX�����'_N]k���>+���c�~�����ӮN�čt� �8�$Fս~j#��wY�K[�9�)�S��O�>�!�D|�4�o��Tx��˓���҉߉C�p�=Q?�01?�E|�~�%_�y&|�w�����;�/Ԍp��x��P��Lz�t0��/��8L�Y{�d���@�f����ǲ�' ��|և{t�c�R:��f��~}��o���=���?�w���C����Q��w�M����}N2R�/]�>�2BTCo?pA�9���T�ČU�_�'�����Hτ#�;�I��r����2��;z�!���k��eVJ��xq8�|��E>��!� 9��/}ł+�
N�k������_�������A�^ $�ey����@p��b�'��ɀԧo?4 <�������q�#:p��3�i�;)�,��aI��JV" ���I��̽��f��#�+/�
�a�X�2yQv� ��ϼeR�6�o��s�W�A�;�QQ[�%���7�����{���?��Oֿ_8�ˬ<�ɳK*���\�q��[?�U5�j�9>x٫���-M��<��bk����,�^���z�����\{��O��N�Jʊ;�v2-%C��@q��4��.	�<��^6�Z�����x⪓������%�5u�w�y��.�V2?�X�tX��W����?���gCǎ��:\w��~�-2�@,��9���3�낆5���	'��3>\ ��?�M^�p��S.�^挂d��̛������~��������Y3}�!�;�k��3H�?��3�(�����L+���/��̌g�?�O��1=�[�+��tU0���>{��C����Kc�˙K���Pk�,���@�PaΤP�A ���	,���G����(�v�/�2v8��%�R�/�����PW_���&ºPUXf���9R����oR08U.C�7���r�S{8�FG>H!O��#��W�W��Ҹp�4><�B���v���'�ãD)���<�g��3P�(����Қ%�s�4;�j�M�%����i\���v3?#F��M�y�K��wߵ��Ա�s)Q�0���0�;b�p�(�Fw�Ěk�c������*�>m�ot���o}��|���Y~A71RJ{Y�}Du"�&}�f�F�p峱���/��2��xf�;��3�A�d4�T�P���?��6�`C_b����3[�y�
�@��;������J�9B�O�����G��БW�W���o���7↾Ҏ���~��M��ŏ�&�����:��{,K�+~��1�X6��P>`� a�NX �b�|'Op�����������|���%f~��\�`����&�`sO�QS����!�	C�Q�1�0��`��J�ٞ#��Jn�-�/�n��v��"�0r�1I�,�d��K�8��{o�t�q�;�O�/�<G�#���(���ǫ���>�:���=��������SaÆ���Y�6�ls�a��}�m�}�����/�s�=]���+��c�GGI�@��W�=Pw�q�]��̖q�6K����D����AE�"��7wF���{��;�ʀy�/�����c?�/�oS�Lu��J>��e��}�|>�O>�T���s�}��q���O�����a����1VF�Do��E4d�3Ϋ���� ~!JV�6�����e<�'�{Yw?���ˮ�n�A�4��(�L3f�r]`�f���b�t��>
nX�������ڪ�(|�pÍ�׿���eU�s�,j�ٳ��������o��ᱜ��`�;��1'?B��/����k�HAOjZ���q�Rx�>�H�0s�}��S�i>�E[� �`И���u�m뭷��l2��/�h���|��W��R�v	[?�<
��qa*>
�_�	3q�wv�u�J��#kl?~����b�clڴ�bt��a����B��W^�G���Pf��`�l���{톛nq�+%��`<q,3L�+V�uH�X�0�&�E��]9I(k|wv����3��4�g�4\����JY�KR�E�^v��s�{ܓ�#}70����RvJv)�	��Qz�%/	��w`�|v�K�k�ب��H��S]eu*����J�ml#��������V�4�֨v�ډ��eG�7���߮_ʉ�`348�zR���u�P�P�����Ϊ���i�?_^�ެ�����{T��(|cC�+;#G���R�$��� o��mg��l�u����U~�veza�w��֐��o3�������9` JK7��,�Y��"�`õl������\���2�v����>��߰�Cm˭6��9܎?�X_N�x�"��4w���+F������:��z���j��u �Gt���ۙ�$�����S���'��G <x�7�K�wI��-�p�_���6��-�џ�'�� �0��HpS�?a4�O\� q�\��a��Oؘ�x',�|�����1��(��t����G���R.�I:�8�#�Yh��9����2�
�XB���-��c���=���2��ʨ(��.��(��ض�b+�~�e��Q\��%�YVW.5�h��O?͍�7��� ~�7�'�u?��) �
b�<p��v�ɧ�ɧ�jw�s����R�P��%��Tk�uְ�շVe�a���B}7���g���W^q������9���1<����1�G�Ha�(����pÆ�0��:d���*��2�ۣG�+���Aـ�e��scv@�~����4l���^J�_��p={˘ ���X_ 8ā��9�K��$��ȅ� h���{��
��" �ٻIK�����϶�n��N����K.uw��	G�A���@8O>����N��.QiV���$r�h�Z�5��h3���������$�=P�A���(�Q_Z�����ٿ�R���}�����8�#�$��S�w����V^�M@����y��Q08F�Q"�0>:'L�f̘1~��'�|l����JB�ȧ�Y����/���R�z�i����v�a;_�����#�mR^[[����J����f��d`Msa������?�<%pf!�gC��S��E��?�0:�`�T��E.��:����#L�Ǵ�'#�lro�o�㥥���r3F}�B�l��N!��ӛ��*�v1W�J� =s,��,�IA͔�%ƛ���&��w֋3���IIb�,mS|ƟUF��ρu�֨�Z�\���W�طR�fV-���k���-��s�����f�F���S�,�/C��.�3S�*5�#	��z���Z�dk��J R_.�m�_�P=K�ښT_�.S.]�Hk���@��I��{b��mSz�ٙ>���̝�1�������Ç;�E�m�(Y���v�i7×�Я�+�{X�h��s� l_�k�'KȓNE�R�ٖ.]hE���:kJq[˶���ȕl��v�O:�7س���/�m���!����$�ա��ꪮ��gd�S�3FD�aiW��=։��]���u��#�N���;�&�b�x���P�8�[9܋�P�h\��@^�����������I��R��'߸����3�2�NPdBݢ?���.i�Gp�)=�e�G0��23�#Kg��PlK�i���=���~Y1�������W;�>��K�)���m'��V�� �ݧ���):Ġ����f�&]҇w���'�4P��1H�^&��		^�X�����߈������^[<��/�e�(��}�I���[�裎�����?�p{��'l�,����j9rZx�qIz��׀�_��@%�Q����v�	'
G;��|��_l��o��r�N�c�+�E���'�1p�/�1K�X�����2t��	����M��݊�J�^�k�Q���u^���Gs�<Mh��(%_d2�1}p�l"���4q��d�gp�X���FA|�Mi �1� ��(C�Z�?1���'Of{��j+�i� �؃~ dRF:}  1q���Ҥcp(�tkioQ��l�M7���>�W�@s�Gc��SO=!�[��b=�s2�֗0������/�~�o� [@���C�jS=��aS��=�ޟ�s-+����@"~h�0p�K�;�7�t�Ut#�3��8�1�j�/@��+�g���ŋ����v7n\w��}$�90NF��b��%o�Ȕ��:k��B���wE�M�,�c�L,��[�`�ļ6��0X��],�c9y͛�Й*¾��^�]O̞|`�\�,����=ʻ۷�M�g�~�7�"�c�dn�e"�*7?|�e�Jp�}b���e����=w�]̽��K��և6aN������2���\�M�f�%q>Wz(�~��T��F�WB�,)��Mz^2�gF�Q�q$@\�5�4�O��^��R�)�L������0d�R6�'N�jhl��̉׮��0��D8uie��*��$da�|rn<�"��;{��TF�d�'~���3E%(3S~���S��#�(���JCÍ@y���ӣ��+�rED�{�ZӚ,?7�z�����ٷ�ei�5~�,Koj�j����v�}7�x�;���؏��;��EE7���@� /�lrSaQ���NRR�r�w�~�O�� �N��.F�9k�uVW��6c��A
fO_�3t�`�����@J�{�<����Km�u��Y$�nF�5je�{�=�O�V-q�����:o���!_zþ�8�K��n����:�\��8E!�p ax��A��D�?�/*���A(���r�tQВ���/i������w���g���G���7�|�Z@�*������Ҍy�τK΃��{4н�����@{�K1�<�4Xj�)tyy9n�^��ջ��C�};;�� iW���f	S V����מ{�:��F�ñǃ�re�3���j��;˙��������N���q?�UK��u� �E�7@�K���s!����	�F�� �,��ڗr����o���=�̳��s��=�K�^y�U{����qR�<���{�?|	��3Ɨ���ֹ�bi5��mC?����F/C��u&����Oy'cL��&����^�Pg��ej�=�����E<��D�ڋ4H>!�0�@�'㕰�~]�b;Aϡm��0p���VR\b�M�l>������V]e�ٜ`��^�+b1��>��a�j�J�`���J�݊$�[�7ޗ�0_��e�Va[Ș�>�����ek���ߣ~�ɖᦲA|��ߋ�D9|����
�<֟���b�7K �d�L6n��$?�;9�qЕĬ���Y?4
���| �+�~����[G[�w���;��Mijl����f�m��E+i��� 9W�/�:�9ӦM[c�̙;��իd�-����<��Ol֬�V]S��%jԨQ�  �����W_�#9a��pJ�tPFO�;��	>��(9r�M6���"r ��+��W�y��a>����8�`M����$X�|��l��)��SO�R!F�`,���G28SY$3�?2��Ğ���$){����(A�ʘ���ٵVڣ�e�HI�ʵ&�kmK#�/{\���PT��u��G��1��K��� 	 �+w�L)�#&[�\������Q^9I�`,����
ό�La%�a9�R�6�O]5'#KV����������\YY9����TJe^H7.�����f�/��
�pG9$� ߐ�8���s�0I���ʸb�#I����<��0����K��R�j���nY��Goۼ�XYa��B�x\#C��U��n[�H �?���]�p�T �eQ^�|��Im���ys��J��X�ZU��
6�tc[e�Ul�m�����۶�n+[u�Q6p���������>�UWee2T&��Y���o���>k/�0b}=���s�K��`O���>�*��;����}��x�K5������?��_{�B0���>(U�=�=�G"����/�0��i���/m�_���A��'gQ����q@���K8�Bwt�ß� {a��J�tCBq����O<o�D��Roʀ?qy&nT���9�z ���<�X>���Q|�h̗�1֍t�C� �rz�w~1�0�H�o�w�e��6�0�eL�
<�����{��W���3�<�a{�> ��ҟ�yե����0�9��w�
?6��[�U.]$c��m���6lK�����Q��Y�:dH0�ה��~�����_b�'M�ec��F��5�ꪍ#�!�w��G<�*]�B�hA�iq1w@�����>5�>���������>����޻�ɽc����ɟ~C�g͜���X��PE�
�Q��ey�o��?���?�<��~���_8ot���`�`�P�`� ������DG��o>:�W�L�|�*��ȃn"$?�wR�?�-/��t�_�=+z�~���͓���Z�Ehz�������(e6q�J���⬽κ���ٓD	8U�H��;4K�|;a��[0���lذ�>������H,ݧ-�{��À�..�\�L[Pk�\��A�-ai[�$3oԕ�E�}���SW�͐�_��ܟX_W����8�{!��W]U���g�e��np�#|Mb�J��Ẕ��Xf6�rŶ�y[$�C-���5�#���غ޺2�6�⭋.�����_<$z�
����ʪ���{�7~��_V^y�ތ.�{�2�渒�p��"�� ~�Yn@�!���� g����a����s�
s*���2��(��={���7־����ջ�c��}����믷�����[w=_*4Zփ=l�z�3J�U$��G$\���ᢐN�][���vc��2��������odu-�v�=��?^�ƺ\�Ҋ�[m��N)��R4exdH�d���Y�p��В�,R��[Nj�:��ˡ��lQy���!�(���i?�*�l�VkL����M�'��A�U�EnZ���^,]c�Z��Ò_҆q�h��9ޝ������D��*}F5����Y�z����i�`	�'.a���j+��M;Ŗ���r �Yz:{���!K
H��l��jϔ���l�-��ق��E�6�W�}��]6��G�gq��5F���;�/�g�w�����P������2����B����t���`H��c��8w�L��˜�K��c���7�D
Jo8��$m��p�'�=���vםw��7d�p��C�E�`���)½;��۳Ͽ`�}�͐rZP�'!\�3��ﰣ͘1˾��<�c+��S�P���?����P�AH����?����P�����w�0,H���tbX��|Yb���<b���<��)$�O�<c������Qf�k�(0(�)�i�8!.<1֍�(CiI��H��.J3�d)'�1
H��b�P�;u(#ߢ��y�7Tf�����~��&�t�M���R�K/��� }pJ��I�P��qx�f�*�Pѳ����:�d��	����T�c�&����j���K�y?��&O�f��W���p����G}�+���q��� &�4��{t߃vxs'�0`Az��d&�'����^Yu@���=t}�>K�⒵?���.�؏���c�^�<⣸�<y�MrM(;��=L�M��~�g��+"b��cH�:F| ���i�0��@|��-@x��_�-���&�?�߆b_��s�q����ب�Wr��٦��T�վ���8�����t�6ȕ��8�Ma}��٘7��+��ؾ��z��vꩧ��q�-7;���j�bA͹Z�~XV�KK��ow�u��V�cɴ�
`�:��蓔���ґ�F�ײ�	C%��>P+#{���w^9r�����i/���P�K�<�1m�M�1�[K��iC����8���Be�:m��bD��u��󺴵'�M�����Z����c������w^Ii�y^�����.�~	0wμ�Ǝ=t֬��|��w�Ǐ���v�)��*���`&�>���r�-����Q�V�nR�0x�l*�P�4q��R����V6nW7�sW丁�;��[=_��^���j�ŗ���_�һaÆ�($KD��y_���Aɋ�;�c�>�r���S����s���q����8V��Z(��\4P��^�`�|)�c/}d������]Ɋ���%��-�R�d$5��*�,��_����#E,yC{�A���ML�w���E��g�X2*6�%W+e�a �h�����Z�I�2E.�TIK��#`Ⱦ޻%�g�X���%a�-}��,1c֒���B-CuRdOm�e,\@� ǈb)�{G+e��@��0�(�w��>�dvP�����&��N�-�E�7_ӯte�#�1�oF��c	�L	Ț�E�p�L1���Qd���&��
W+Ň)��ժK����?� O�v����@:Y��靲#�"m��RhZ�Fa�D��gF
�O��}zJ9��q��%���$�E��A�(|���W^}ŗ+�u�Y.؁W��q����λةg�f%e�V�4�/�� %�ǟ|bO=��=��c2�fJ�8�V_}U���	_�~$���h���/���N�G�?�<��R�5A�/�� ����u�Bϱ� ~y��>��2���BB<��q�-�� 3 �����z᝴0
	E�!}�� a����@��͈p��,�b6��S��Gy)#gx�(��{�q���WحH�����/Pq�����'~��xN���������R��K�0;T/\�XYY������G��߳��}���f͚�e�Q���u�4�}Dk}p������3�nI�5r���h�ߪs'��p �2h��Q�d@�dԽ��V���K��UF�1�?���2�XfV R 7���$�g�Sl{�E�:�c
?��0z�|�A�y���bāwh�/ ��iw���.��v�G��s�6��t+.se�˩0;<�tB�=�D�d�H3�"x:r��M#3�O�i+�N��w�c:�?B|�߁00^�l�d�*��b��r�m�����"���}��Ǣ�ul�-6����<{���Q�ǟp�/'�G�C��N�Ϙ9�z����99�ִ؛o�mʹMGodC�J��n��l��h���'QW.�8`��H�N�6��<�L{ᅗ$�� @��M���
ϡ���pW���/ClO�w�5�#�a��Ҿ��v�]t�v��O�3N?MzI���>;ї�$+�=�Y����i��l���v�eW��ѣ��� � �9_��������2��2tğ�-����z��j<昣n?���_V�}nHu�ҡ����_|;qb�o���x	�㮾��w�~�;�H����Է:)L����j=�\�y��E\ȉ���AP��,�@�t":-�5�C�[S�|ci]�=}?F}Cu�b��z��7�h#[w��l�ر~�)����sO[g�5-S������;�T�A��Df�C.2��] �����|��F��>�d���s/�m��=�-�kE�[U����k�>�Y_#˥͊
{�$�z	O�8��aM5� !�ꥣ�5�Z�t�L��WSKZ��\k�R_�Q�A#ǚtqJ�G�J%S�R���(m_NCTI8墹�	��F��η��B�i-�V �(��՚�+Y�y��_dm�R���$���Q��T~fפ��1����Ho,�khQ��ZQ~��~X~��a�סh)�v[�jaV(������$yת�/�O���&:�U���C���m˳��v�^2�/�%����Ysk����h�S>���Z�"��2+��|�YgّGA��]u�uv�I'Y�������3�G\~��HYy��4�:��bf|8�/ZG�GEO��|?��W��|�Ͷ�6۩o-���;Ϯ��V޳�8 e��~�-�Ϙ>��:	G��ӥ�J�yV����g�����9�XW��o����׆��7Π�sf�M�c��T�=�����?'5��e��QW� >���`�3V<3:g�8q�7����S��B�(���4�?�g���ₒ�!²%�,)'��4��̔��M������)���Ñ7N��e��C�1&�o���n�ܘCnG�����bP��@3�0���EP�P�G\��*��(7xf�&y���%�ܝEY�����l3��ۭ_���٧���'����i���2hQ���֚k٢ŋ��{��a��U���S�r�`&35_������X���ԅ��-��2��J�b�_�.�1iS_�E���"�����/��c��w�O �=�>.����7�'iɢy��)��Z�h�iH�.���w1��!�/�Ov�Е_*�$,Kh�vc5�R��4;�����������`)5���h��v�/�g	��믟�;��0k����?�s���������,�&ݷ�~���XcM�P[aA�-�\,]���{��x�w�}�](åZF:
�=���1���,�%�n���>�;��C|��1�f�>��z�av��/�C;$��5̛�D��~��|��͏����hg�q��0�?��IP��Cք}M�u��Guԝ�{��e�e+������|��}&O�|���Q�]vY�7ߴ��9Ʈ��Jg01ܹ�k�]zi`��hi�D�L�S��
&�L��)0 �aΨ�����"h�aF�W^e�(�����Zwݵ�@F�mw�mǪ���]f8`
1mO?�9���3τ�b�=Ǖ�>
�<�����:>b}�CO�ՏfEe��k��u���\��^�x�͚1ٗj��n��q�p����t�4�m�Y��l)��g��R���Y_-3'�r�^�FM��yKPNi��\0�<)D�m��P�ࣛ�2b

�,C�[5q#I捵�I�$o��M!�-�WF�j�6���Ϸ��rk�VaM���*G�,��69J�*#��βs��D���&��"#;�M���	2���X/.�P�(�������5KYF�8���++��@g֫���V��eHi-���ɴW]���ko����6�����l�W�X��)�ֶۭ��Y���4T�FF�Q��\�X��ƛ��c���na)� e�9����A���Ѕ^�S��X�Qyf0��Yܛ�o�,����t�M�d.��Ǽ-���t]�h��>�QH���)'�u��ݕ�q�E��}������駟�;���Y{�/eB����}r(#�生��ue328�G8�$�E��4�x }��/�I3�A8���}vEm
��~lW�&v'�w�E>Q!��"�W���Y��Ǎ^Ҙ3g�ʲ��u�q ���(S���{YW�&M�,÷����O8躱�Q�ߞ�����m�����| ƨ<�z�K���t0�X:޾��+�v�����n?�i~���~j!'��6 ,��rou�Q�K���h2
�_X�x����d�M�|�����{��|�����Ϊ+�z3ȑ�)ޕW���wC������%��e�(�Ol�dp�.��]�D���������6��%��3N��v#^"��-�O��Gt��
�'���-~
��`�h��]K+����QGm��z���D�0��o���~��m͵״{��z����CMm�]~���#�I�Gy���^~��Ez�����w�������O���p@
0k�lGw����Y�ŋ�7���N��ю6q��{�QyKm��ʄo&H���?���^=�1 3��S��V��֫O�-^2��͟k�5M���|(G�7ַ��ǝ`�����?�V[u5˒ld�Z��?1�a�9կ��|�v�i�y�+h��ŧ:[�%��N�Y[[]�QGޅ�Խ���D���e�r�����?���W_+�{�5�\S��/ءbNz�0�;k��z뭄2�&A�l��ft�
׹[���CGe�F���x�TP�:�Р40"�R*����N��H0Gg�)�x�mv��b��+�����p��s&���
���<bz���W=��������«o��`�}Z�!+�R�nb�}��S��v�B+-���&"L�����o�mV9�.6�6f)_Y0����P��r�wQ�5H�i���Z���hwks�[A��n�-MiVt+t#��mJ֚��:q��6)�JI��.CId�e�JQ�4��V��~����[�и��6vf�M���*#(3M�cKۤ<ä1�3s�Z�&�	ޕ~sks�MvV��˒�Γ���ʻU�Z�0�7�'�����Ub*#?�曔u��V��o�2��͘dMՋl@�6�o+���p��������+۱{mh�L֬W�BX䳖�]q��~�iֽGW��3e���������?.�
.�M2��c~~���i����J�ڈFX� Yn \c�8�p������G(���^h�=��=��S��X�>}ϔ��(7�� 8g���jL1���D�)K��w~�3@	��N��ݣ�����~�"9-7�D���$7�}Zj�1}Zx��eօ���$���9%�b|�v�N�:���y�(�H�4(������g�#�p�f<K�h#Ҡ^qf�8��b������$~����~��w�Ÿq����ۭ����7�zs��FѠg	��Lws�L^��q�<��,y#���G�q�1š8��;3�,�",�I܀G��ټ���*�b;����I���+|�o��~)��=�G,�����_�(��-:�G��?�%��%w���"M6��@L;by�]2$�-���U����Cڕ�b `�p�|�u����_��1��Q�ɀg���C��;��X��9P �f̘a���?m��ڰ#�~���g�p��2s����:�a��{pG�6�l�m]rgˑiN�&l�J��d��⇥��6h���ꪫ�Cw�>����7�_o��Fv�A��ћ��s�>�=��۾��k��2+���o��e�-M�nz�]tх��[`8�����D��8���3򗿜m���o��c�=��8��h�P�e$F%H���M͍��q�g���{t��@��e)r��a�w����㏏�bṱ��Z�����aG��B�saI���+��M����@���s���Ȍ�#s�R!��a��oL�!�)J0[��e���;��%v�ŀ���(�����s&?$T��]҅a�L��TW\y���V�1�R~�+(-���a�kmIu��w�f݋e����P�9�
�"#Ie�n�, #Tl)�߯#�%G
a.Z�D� a�Nʿ�C��t1�,i��Q�P�Q�0fJqi&]��)���巴V���[�ozM�_(��³³�c��9V �}�A�������oM���*{�ny�'�Ii*O�ڭ$?W
��?qo%ho�GJf{�l/
�,� ^������5h���يр��B}�cT���dVJDfS����Up�܅�TWo�ʋ�L�'S�}�-�1��m�#��a��6>����_��}�r%;8�[tИ�6�����o���a�(߼G�-�{�d���Ӧ��.����'��h�/ �����ɓ�G^(��N:�o���gԯK�WE���!��Gm��2��&�:�4Qԩ��u�EE���0�?�:(�oԅp8� ݈�ׄ�l�ځ����F�1}����?u'<�Sv�%�a�N]�'ҧ\�= ������~c����~�%,|��,'d	Y]C��C��P&�&��h��g�#b�X���!i��n��!�n�\}��\{��Wl��¦xx$��7�|�Oc�'��ŊY �A��9�D�l@g�W��$�}����N#ڦ^|��HY)�����>@ ��:�x� ��Q�dHއ!�1B����i���L��ԗ��7m.��i��b[&C�;��R��=��@|��1~W���0BK8�Suf/�O���[1���,)���I�3��=�ӧ�@��U�	:f��~��5T���eݽ�K7Y����n����3��$�@��+�(�����窊p�3y�~ؿH�b�����l��v�o�]q����v�q���	'��E>���-�={I�ը���p�`(:Ufz��qڙv�W����}>�`��ys�O]v��v�a�ؓO?�����x��R�8$}$��L�}q��U�rȵg�~��e%eV�/����_�o'N0nܸߋiv�M7u{����c���/��� q�#!�q���X�O�ؽS	#�3�����U9RF��y���/���
�ߗ�B7���Я��߷����:~�S����H�f[	�̬<[�d��.c���Z�R�f��.�Q`�U`o�G�$d�`�4Y���j��b��TXUe��-C,O����� ����6�1}V���C���(��C�:s��p�M��ܢBkW�4W��)��(C��a,����U�
��_��J�*��X۔�f[�8�9*c�[Շ��2d4��ڼye�d��fA�kk��Wo+.���#��B�/�b�� ��M)U
R-�m�`=*�Ìr3z���'�H�t]�o�źcYT��+FQSc��t+��G���7�&O�oo�9ƺ�v�]�m�(�zF���O9��BX�����n��X�
:e��-4�/~ɀ*���d:J��N�(����Q�(@���=� £p��B^��C�`��Ϸ�6���|�-?j6���5@Z�%��H̍X�F�`�,i�i@���R����:�@r{�����Q�&��
K���,z���݃�OyIG)/��b��� �9ΓBzY̌a(	�Oe�R�#�2C�8Ҧ~�2b�qI��	n�O�Ƕ"O����6�|�hC��o�7�đ8a�ugv`Z���(!O�Iœ���O;�J���'���>�yc<uq�6��_}�5)q�~�e�|'-�@��3{0(x�}�/�;��.q4#|\��XҤ�aa�/�Nڤ���	�İ�&;���?�
1���x1N��;����X߈;�=��	.��?Bj�]8K��%C,��~J*���`�RF��BK�p)�b2�H�<�vgi4i���џ�)���"�Bz�ʋ�Y�	f�
x�xa�'��0K���/����ꂬcP "q��v�l�8�����s����kj��1�m]�w���ڞ{�e�uM��jk�Қ*�:�k��|�ć��j�s����{�y�Q��#�)�ޯ��*+t�H_���[l����_~�9�P�?�ϚŶ�B�l1�����ru�Q�t�I�IY��5X�5��φN�0�T1�o��ւg�~��Pg�t�
	h�.H�Ů�o*�^@"͙���������K.�?��>�	�M@��� 9�	�Q�'C��/̝_�@�4�%$�����c��F;�@3A�넘6�8�^r~����!�A2�$�xV��.�e楾�ο�pJ��=�F�>��f�������T�YV6w.�GD�UvH�	�R6cK@���[%'U/�fN���R�14dp�Y��pʝe%ݭUefd����O;KoW~2���:d��=�!Ų.NJ���Au

?�����������=S�XJ���_`Ç�ee�_1s�\�#�/;'�����A'#����|W�YN����k��o���>��c��Az�p�x�BC{����-~��bz����	�XT��!���
���V���H$��ŗ^j���{�='2��%C|#�I����B�Q��L��� ��:S��%jaY]L㊴x&eF1
��i\�ܣ�S�ph�ˁ�C\FL�����KB�N^���C:(!M�+��=#_ыZ@aC=(_����a�L�6�Ǝ���A����?�1�R#e�����im����C�bX����q��=,���|��|�~;��n��v6t�P�'� o@��3|���ɲG~�9��[�^��]�?y�ު�������@����	� ���]��q�"@Y)�
��8��q�H�4b:(�|'�}�g��_§�<�ˁ�t����K��7�zS���S����tS�$8I�ѿ��-$T4��,~K��v�>�N¬�S~V���"!,��-�!���@L�8��I�pN7	]�7h�6�𔠧D�?�$��/o��v�q�m'�_y�]���%O�m��9�[ڥ�^��A?�p���>�ti����}��x�� ��֛lݵ�����%G�l��J��o��^zֆ����q�.���o����w/{���Ï�I�SZ�8Z�@���1;'�RF�e��r��E��+�~�JW��yｕ�L�rzII�od �<����b���UW]���C�D�!tQx�����1�ѣ�( 0.NDb��g��D��B�a����&0��<�!�K�7����k}��w�>�������J��-:�w&~(e�C�y��e(�hI����(�> ],��Ah(h(�ꚦr{\��#UNg�u�/
,������uA�OE�]�dg�t!�LLZ
���8(�8@�q��R���}k���B)I�o��
z�6q��=�g�Y�\{K�+��(���?k�30e$�L��`�]@K$��e�Jϝ��h˿%��7~��K�bE�%��)7�X�.k��3���&G�h����@�t�	���Y��=*���b@� 4G��˃�h����.��
y�����O���e%>~(�5UUv��h����i`6�����!�9'+�S�#�1���8�G-���c� yп�9��X\s�}m�[�5.�'�%�q�Wh�0��LmE�c;2�M��.���z��y�];�3�KY�N��4�mذ��S�UV�%��C�Ӻ���K�a�=\�t� E���1�C?4�
�?�4�QNҠ�~�G9���	��
K�EX\�������	�U��0?�]���U/��E�Q.=G��Nٓ��
��v��ĉi��a�؂�v�0k��{tΌ&�����5wԋ81\�ӈ��ZܿD�!9?�C���~H�U	�3���҇lםwt��]dW_u�����fϙi�[�袿[~A�}<�S�s�}�ri�:����m��&v�M7W(���Q$]g���v���o�bCu�
��l!O���z���7���|Ď�0��։#JM��q��F��m-�G}���ß�,+-���~�(y�b�?\y��is�[�G7�s�KI`6t���a"�9���)/7����P*����5�P B�5�|�5YJ�|ȃ�s����3aD��ƙ��� �8��˥,Q2�(2�����{�~R� ��iE�ˊ��i-A�7��YɃM��2�`b�!U7�'�G>2�2���2�`��ýA&<�w�&!�ȟ��H������`�N�w�T�Z�Ia8⻩�яT:|��3��fˀ����`�`��>-��J�ٲŴ3U�&�U� CMF-�A͊��i�#��j�*O�����P'6��4)�,�H
���J3(*����
D��S=�k�ѳ\�g�pܳ窥��:�9=<��2�H@�
���O�='�a,����?�Nc$e�QFA�D��2G�dH���w�x�G�K��W/��ǲ���i���z�%��Q*/��v���z��ֻW�S+��A(,�I�63��������;��\��c7�w,���6,sc �B���Q���o�Î9�)f�~!%�@�C�T�YK��L|�x��y��W��~g�7�Z�yx:3X��G�r���ih�@��IߏQH�oN�	�����t�׏���Q����u���.��g�z&ljک�� Nj:�.�)��Kqj՗��g.1���	�\����_��������E�DK���}��Ƒ���܏���<�o�BN&%���@b
�AO��v݉��v���/��z���3�=� ��ҋ\~����^���E�m�����}�j�[��}}yU�نv�aY��F;��C��W^��F��1kP~y���[� ��o��N;�d���u�zz"F蓝�2�V[WS{���z޹�]Խl�E��+I}�B��q�V�:u�9�{^}�U��ƍ�#F���&�f���<����蠡�:sr����Z��ѹC$P.��%0R�rF��P`�� X�Nx��5��$y����I��a(GpR�t�%#��#B`^bޜ� ��q�d��2�7)�zQ����p��ZBC�@@p+�4�����A!	���!�6��1B�b���a6r���se��r<%í�eP�B�����2.8}+��ղ،��\CuKF�L�F���@a���a���.��o��%�������&�pFQP����QGU��{�18>0�8���1}\8�!�M�)zܡA����M���zZz'=O�<} ���9��h�=�z*��"���f:�A4T>	�a��7�(w�o�K�z���{rV_}_JE?�~8�����i�5� t���$3v�}����!��\����.�˦��4�Fq�)���3�l����8ʍ�KU=-++�0��5��eY,�����A�?�\I�4N^�^�g�%�r�_�ߛ��|�0��}��<���y'�p�u����-�:�-�7�������5���=����t�h[ݵ ���!<� ]�WTo6{_p�v啗o�޶ 8g���N�T9 �|#ԙ2�����pG8��P��G��eT�_�D�e@~��G�cH?G�*Cߎ��a�'�X�d ���{��b^8��4�uO ���y�;.�=!�;b���@j�+���TY�B�3�>�މ�HF��ヲ��B���D=���%d��/�78�v�6��3KK�ȓ�	?�3�f`i���~�{�v�q;����w���-7;�����c�v���>��#�GReU��������gO�9sfJ�q���o�ު����C��g�~�V^��^L����ɓ�?�x�Mvء��8�,�o�vǳ��S'��7�yCmmu�1�s�9g�s�C�w :_� �0a�J�}�ݹ555{�x��v>d�P?�5(a�Gd<Ҹ��*g@	��G��ľ���L|�#K��Sp�	�a�������s"�Thm#5���&�-(�kz�5�p��_�e� .�F
��~���~���~\P?x���3~�����y)��UJ%�G��9�H,��2�bۤ����o��1Nt���M;w�Nl�7�������ŋYS#ʲ��1��"���1���d�#$� ˬ��e?X쓔�� �8�ad�¢\�e���
O�x�c��VTp�#*��M5}��f!�w���������M`�Ũ#7ȡC)(���oh�p�t�7y����-3��p|�t�2J|FRe �ߣ%���/���M���g݊�1��<�-Y��/�ᐉ����m�}/��SUUm�L�����=(mD�x^��0������_tQ^�P��,��!^2��^�CuJ�\Q��L>??'NW�ZO�ߕ�ρ�dΩ5�
��%�p�P�%�"�}�!���o��ǽ��6[yܛo���9�l��>���rg�p)+)�W_Ï/�7g��AhIT�h�@G����v��7���<��z�M׳�s
�q���s�Xmu�H��;��{�N� x1�b�=�eZ��k���jjj�9��S/9�̳�_��~
[�A��oV�8q�_1�n���4�:2l�w¸�"
.Od>,���o�{2�N��_2p1=b�H�4�b�Z�i	��|�7�����+��8���O���b:?T.|J�SK�\�����Mv�E�����.���w�E9Fy'TN�BqW�e򎳱�cD�\#ġu�	BZ �ڈFxIc�%����w7,qR��q1����ׯ�f�е�o/(�Ee�|)3��1ᗀ���2fܨ7���t���Q�S�_P�e�%�f@�a�uW�
�a~
��nL�r�\8��2��Z��0˾u]�	È�׍h���c���S����^ϔx����w�2�T�w��[28_J�\��خ�Oq��#�裏�qr����a�g̲�ƌ]��@����m�5V��͘wޱ}���)�\kmZ���[��a�dhK�,�����>��4d��m�"]c��n��������O>m�z�o-`���򫗨^ɭ�jkk������3N�ۙg�ySQA��D����ˬ��� i�	&�/���${G��O߾��at�Ύ�OXR6��ac��� ϑI%3�T�e��2* ���	`q��H�BZ0�'�QV�}/����d |r��C��oAWuH��υԴv��x1�屢�	i��4�C��&��Cu�?:�"�B�1��t U@��U�`c�MX��9K�?B6��P��쎄t�@/1^8F��f����q7���J�]�q ��?�Ĵ�%>ߘ�i��b˶�C���#|�	£��y+�R�4�#�3����8��0�8�����~�̾lT�ϗ�;��gT1.�i�KF�Y�{2c~��z��ж	�R~8��X�d�/b�RӉy�쀈3��������$�#���~��CWu"ʂ��b2Zω��7e�L˃��Zx=S��֩�s��w�2�T�w��O2D�J�q�K��W:�5N<�$;xס�f�{�Nk�
���#v��qu��2��Ra'H��6�y��𻉓ݘ��/l���^vh�_�p�~���m��n�f_�����#�r�=H��WOQ��[C?��nKks����O?���s�kV�/���W��;���o-�i��lӧO7.eemyaF�L':6֣P�Ê)%���q1^W��d���t��L�Syőmd?����~~J��� .e����:����v�����)	w?Rc�tR�&��+��_��J��yy��*]�i�DŚ���t�#���g��������`JT&�i��LzGY'<�o߹$�x�=�ؿ���� rя8�/ �03F�|a�2�X�C}�hg�ǲļ85��d�?�54e���$���D�&�a ����ݿ)Lǈ1+�c޴�Ƿ�W|&Lr����T��;��t�Kvgˆ�u��@j��S҈�Bޱ�r����of �H���KH�A���+�ּ+\�⪫0��U��C�c&i�~�?w�q����m�)rSm��6g�<����;ﲯ��ڏ�>|�ߣ/�gFh��L�:զM�iO=�����Ns���/)�6��ǝc��{ڳ�>�G�C���H�^��a'N�gY{M�o��˛n����A�&�����S�
��_~��'�|r�:�n���oXE�>��&����͐t��|蜝�m��H�#N����)3HRQO]��W���wv@���¡ 0�6��BL7Bj~�r)�<]����߅嗘��q �Ժ�i�矂��࿉�W{&�K~�8�C3b~|�$���QqGy�1Ͱ�3}\̓���i&?1���&�,��H-3�����2�o@g�eˇr� �y�ACt��^	�%�.KI7�'����/�'�˃��� �G�y���f�5�����/��} ��j��.@��u��E���v�}��Ϯ��z;v�+ʑ��|)i��$�U��Ӊ�R��_����W���_���!��?����&p� �5`h���o\�$�4�U��$Tfk0h�5ǈ�2���L2xxf z�:&��)\짤�3�����⎲��~(��L\��ۉ�'B��yd�-��o�~̑��3';'qA�
���O�BW�ԩ��9��t���)5bM�rnE�P_���u���st�WH͗$�J��뺸����V�V�I�A*m��b~�����8{���p��o��'ǉ��=BL#򢮀bp�_�v���Wi�r�$�\�_r��o1]\�_e������L'>/&��i�����d����s���K�����GH}�wCr�8��aVN�͜5˞�y�9s�+��q"��~�<V�������FX�l�ĉ~�FG�Ϟ=����������{��U\w�g{�UYu�zA�$	D z�q	��`pM'�{��؉;��q�`���]�#	��{���^����j���7�����y�>��=s��is�̆�mӆ~��C�|5��nR1�2�s�=��B>��wV��"�y�fc�'M���w4��YP�I�m��2�{W��A��@:�J^^^��@#�))���)�(�8𴵥=�f��{�J��������<���p�����[�o��n��J��н"�c�����\�����������=���+��}�^Nu�O��m�|��{O���������tC�YN�n�	t��P��?��+�(���NsԞ4y�{z�;�t�C�.aL�j�z���gy�����wVc6L�)�8Ȇ�(K��5�/V%;������ûп��������յ�!�lp���'G)p/b	�MJNjOKKm���k ���$Ao9���B�&XkCC��iP>��{������^�_���^�C��ؗ�w�������D��$������>i'*=���=��h3��������흵��`�t�%�k����ҳ�S��r�������u��.��w�F����wB����j׼�ӵ��s�S!����F>m���q\�εV5.Ӭ8��֜0��|'�'�@|��i/�޽F^G��$Qy.�Q���%�ݝ�l�ͧ`oOJJ��q���+��iV4�49��N۬��^��܃E��{�����}��}A�<�[DX�!����*�I���#�!N��#�Ǖ��	c�C
�o��
0����Ρ��H|/�φ*��QU+^i�T�;�'�w^׋�����o[���R�������\���z�k�?_�?=j(����M�B��8�zJ�Ѻ�y���nq��'�R%@6��w_�u)3�z��b�Kʩ���w��o��ʵ���v�N�V��� �7��Ʃ�R&�7�!T��}aq�y�uO��'�����+�x��s����T��?U�[�{����� �ڣv�M�u������8�G�	x�/(�{=e��?W�}=q��z֮ҝ�v/]39T�n��M�xש�޳�|��_P�܉�結d�k]5�i�5<�o�Qފ�PN~tE�]����M͖��j�z�{�}u�ޗ ��i0���c�
5������)��$�b�'5�(�7�U��L�<;��v�/���o����~�wʟ���Z������[���'�S��o��V��!{o��d<ߑ�3�\�on���h(Q�<1��S����gC"��%����s|��R������.jp�.u'�n�=����)���rM�$M�dM���1I�YB��cR�2�7�kb�\��=�s|?�{�䩼E	���M�H����`(%��P1�R�Jd�r�R�0�����OV�2�d$���v��1�vI�5��x[	��b��`�D�����Y��,]��_`|��Ӱ,O��;޸�v�3��Px�;q���͍�'�]w����#���:�
�p��>%���:��:��>}��[�BR������'ަx1�CM�Z�%h�q�)��C;�x�X1��Hs���'|Tƿ{��1�wa��w��[O�����1Э��:���Q�6�6�!��W7V��v�]�?��\vzD�'a�xxO��+�#�h�3q����;��R��DU�'W�?���x�թ�OU�鋮w)��KxC���8=���s�kܩ��v����P'��B�_P�C�׷����x�J�{��-U�y?���� �<=��٭�,����g��ڣ���^Ou�g���N��{�wy�*h���L/{Br��O�z{���Y�`Y�6��4��,`x�5�j�O�����ۥ���C�
oa^���K�{�AGtA)�T�ܡ�����k�7|�.��翞�'�y&^�^{��G��>���==��yO��(���\{�`t��n<������]��p���^D7�4�/��K��v7~w��i����ȯ�\���;��'��%�p���ݠ�-����-�WaLR�\T�=k�*����DI��d	��. �:ѻמ%^�����R�`���4�� F7�R�]ꍸ���'�J[^�X�<,�"�&I'�C����(%����50���;�'ݕ-��A�;��x_��F{�r����m=�bFh�?U)�]�x?f՞������� �UU��</cS����d�X�V�T�0�-~k�����F�'}��W��O�
%*n��m�n����ƨ'|���߳r�B�a�B��q��e�{]�Aӽ#�﬚�C�bZz�t�f�E�+���<QO2V:�����'�`pj�$%C��FԠ�+*%f��x�^OUh�{�o]�{���GC�������*�����O�;��~��*=�������	��jT�O����/��SW��z�y;�O��g��S�O���酂�?C9�ʉ�z���P�ڳB��m���o�����UFRZZ���$ݣ��l��	�A575XSS�������U�j(0�?�K{o�'�;MP�k�j��=Ǣg�S��j펻�J�x����==����ygW�~����T��so����o�S��6g�[�^�Y�֞����,�-��;`�YѤJHOOO�GA!�lM͍�����xQMJf2jb2�bЉ�K�����s��D� e)���^���6k�o���F������ki�Ҧ[B�fg �@؝>Ii��Nz�K�w�HN<�=��3՟gD�߉��]]FQ�텔��L+%.��H��'x��\�ʚ��U_	;Qa~> ��X���a5]��=���{D���}|&���O��俧�{�u������;�2l;����O|�o'�X)�L�Ƅ '0�a}��F(�����nW�Z�?U㽔`�w)��2�=�`�t���I%���4�~$I)K��R�N���N���ƚn��{��S���RS1�y/U�F�0h��+zdx���ݽF�t�M����,��yA%��k����l�!�0��.�{�<�����f��?����J?N���M��X���^O�������'�����z���r�O��d�ƸB+𥮹����ڳ��K���������Oxz��V�7y9�x���w>5/S�R�2��i'�ħ�$�Q�*U�������\��
�:n��o�g`����v�!�v*��\#��\���)0�M��ΩƦ�=��߯�b�G�h�����/)�zO��R�{�T0���$~�����E�)|�7���������"�����w�N�RQQQ��k��ۮ]��x�l�ʕ����Ɇ׬Ս &#��ΐ�J�_������H������5Է[K�mW�����i��X���Ԛ=�
�%�Y���]�I��C�"��B��{[D�(��P=Jd:Q8tXl3��{�+����B��M�9��4�F���3#C;?���;�$�{�C�#z��oA9��;�ՙ�z»	у'�N����Ca�h�g	�S�O���߄Q���_�Ȝ��cu5����"%�0�$9tE�[��"��h���FH���8�i�%|F�&��0��u���R�7ǲ{��.<���X"�Sy}�χg»��wr�����(袐�iW�<T���N���<U;/���L���F��H�������i�g� V�zo���'�?����.χ��I�(����� g�1�P��IEt�oQA�����܏����.��-��Qh�g9յ��ϵ����_
��E}�Ac���[:?cὴ�}�3��X�-�ěx6�q(8���|qc��pG��'#���C�x���L|�6�\�>'{���X�n�^�_�o~km	2'%9���ҽ@������4椮�_��{��E�p񎞅nrg�mឮ��'pD����m�¼�Yh������C�ڽ�����/x_O��|E���w/��˭?_z>�>Q��~�}���]����/(���|G1^ʶ����6���?��]���&'&�=�z�iQ��T�[����;w��jժ=t�Ьy����ի��! ��ΰ��A�1|AYc�#�N�{`h�ͽ��Q���&�%�{Xu����>E�6�t0i)�,�Y�f���#��G�����gEEE���v���B!I��/v����aia�R�P�V	��fV8�D$T�@j�R�i(DF��;Ϸ�5�߆�4oO��b(r�լ�7�;I��G��'O��,���׻qTy����_]IIM��e%&*	���i���`f���p�dIP���
^�ʪJ��)6�=I�'�#�0VA�y���J������ ��a�`�����D������ ��$�N�*h����۷[��r���R�a�Y��^��(�����ߺb�yg�-hP��#�S�7-2~}eK�{��ʃz���f�;���}q8�͘��M��x7����>�Jh�~�Wh�g�x�t6��
c�xpow:Lh-���C��tC��t���lx.�>�����8�zh����6Jk�Z��w� �����wnn��WGi��W[jQ��N����,���N8T�!*�݋�K�q�bp t=�G���˰��/}Hռbu���肱l�>�rM/�|m�.�B��6o���뱝xO���x��ߔ؟�v�v(�9|~� �u�O�q����~��S��	�����W��*>C��R��ͳ��pF��ü��
1��~o�_���~h�O���
�\�m���B��XWb�»"�"nb�~~�=�0qͯ��u�E�N$��0;^�z�)φ�i݇� �j�]p��mz}�sŕ�\�Cҡ�{����q'4�k��C{�������|�S���Z�G|_�Nᾞ�#^��o�S�iu�Sa9��A��L�dm�)Sc��=�a��'މ�Ɔ߀������w�Ả��?ڋ}�������c���w�9K��mt�Kl���}��[��3�Dx�3�Fg^��(|���7KKQ,� ���<x@�G��o|��|�Ώ=���z�@�-�m9�rz��zY�v�ԭ[�����?��O���_gZ��|�yF;���f���&V��=��Ob&�*�':�pF[W[VV���K��؝w�Us����n5��v�W�����w�{�^x�E+�["_ko���9r��I�"�����{��P�e5[��oa�D�L2(I|�0"~k�w�4�"6�{3:9&���Ld~�dıB�!pK?Ç��3gڥ�^*�t���?�];�Z������a+?r�[�L����K����P���_G{�:ҊK�l��VSuL��?��s�	��Imt^�u�K�u�;^��6�t���n)6��WI�� c�Mc���nyR���_M�u��.E�|9�t�]�z�+=���C��,�P�(��}3KM���ņ�6I�2?` *��(V�?�[J�+_�OJ�'��ċ�QG|�����ɥ'�����whz�Z�}2\�' Jc��څ��!,s�D6`���7�7��>����x��:&Ù��О}]en���ūM�I��Mq%H��"�Q����c��aS��t�a͵�@�p����:�S��ߙK4��{�RF~�>����{x>Uth�f�R���'���^)Q9�C+��6�=�6�n���P���Y�����c�wڠ��$U�H�wZY��ߡa�����fQ��^P���;np6��ֱ!��>3�y��|�a���7���I�5{��s�u��?�_�/�ɂ��cHGTx/�bpD\��d���'�q��f� �?Z��ٹj�����gT�����&4��W�Q��2Ca~�J�"�ze�x	����ZzF��D#���{"T�i�L��K�/���:��x����..c<�l��$�[����8����߂�ǉp��w�����Q"����:��7�#}����{<����+��ݛQ{�Dh��qʑ�"�ڀv�����?�'~�~�v0�b�~o4��I����}�����q���w��^����8�b����~�_�*/��w��wR�=�����=\7�r�/}8����l8��k=zĎ;R���|��w}�G��`��/=髷�/��۷Oݸq���?>�����mڴ�>z�vÍ7�dC�2�)x����]Qil�+�b��5~�4'Ms�8'L����UUU�X�$6���L�>�Ŗ��ǌcs.�����k2����J_E1b��3{���[�UT�;�!/�C�8���ͱ�cǊ1$��{e��َ;m���V��Z�W[gUR������?����!WRR�U��;<���q�L��/�a��V�Zm+V���¤Q����J�4i�=��c�����������<xA���WTG�UΐY�8�F��'̺��Ib8��ikk^��9�N�}�w�޽����HB<�?ug���Cm'��&}!4����-m-�$8H��,9SS-\I8c��j����#�M����V�Z-7'�R5�I�)XЍ���%
J(3���^��{Q*��a�8���)VϪ�T�4Y}#J�ER��=s���]Ju���^*C�H4�AGߩڦ������쀓V�uu��N؂�
�D�0���{Y�o��3!��q@�@ɥO�j�ߧ��
p���hZL�A1�纏W[	K���?(��u5mО�g����E�V^ϐ	*$:������w��;���,\�*��Pj���ʭ����^/��ǋ�����.Ä��� ��������	�㰡�7
&m���`p8:�����g�-����Ti?�?)�F�r�'p�q�0�7c�3�Bߺ��U�v
=Fm		��Y���<m�+cE!a@��4_�^TX��C�j��.p
��#���+}��Cu�R�o�bc�xi�h\3bл��l*<�q�7�Fz��(���yN��}�0����\�ގ��6�-���@Yx7�N����Gh��i<��8Qy�II���ߎ�D�8q����7W����hkn�(`����?��y���#��?(/��=��@P"�%C�o)���Th�v��>�AuI_x_���}R����_��"<���p���: ?]��)��-��A/��i@b��ɽ�����3���v��.Ń|"�/
|*�$סƙ�>���+:i�[����-���Jl[�� ���R�kqnA��3;O�=��yƯ;u�3�O�>�A�0��%�|�H�1[�[�~�[���'?q��!v��9���t)R�',[��k׮�����Px��m�������u�
�d͚5��� 5��R�Q����4n�8_ia����!�޳t˔����s�Y�#��x���#8��Y
�8tȶn�ak׭����PUx'0�9t�P9j���8}�>�%|�>RwWUV��ـ~}�@�
!$���!%����C����}SQQ�mٲ�#�#�X]Sgk6�&�����uz����BmM��'�ZY�2t�p6�F������)ŕ���V	�/m�B!�wF�~$vSzP���q���C�j��bTV����e�n�:������h/V�ee�ب�#��b	�D+,�s^�,8t����0�o��~�Uİ���gVV8a��/19ECEc���MR�j���cG���=�e ���e���%aI�QNn�6�f�?�&��>��P�7���O����~=["�5�==��A�s���m׮�m�V�4v��a����2.<���!�(�A��ȑ#mذa�`u)5%ս�)	2z���.*m1�|2W��LjEC�33�5�u�@ ��}���*���7��pg����=%%<|����e:ɩ�<�'��A�������w1�q�v����O{g�{~�y��8>4���Ç[y���j���16�	} Oi�@+�ϱ��l�V�N���d5��	�$����ը��~ƙ�d���ZUU��x���G:�w�����AQ't,��~~|,��	�N�#x��w _X�����$��N�f�.�Vuf�|A{����N�v��O��o��^r�%n�C����P�ZD3�/����Sxo|?��;ΪO��8�|Mu����PV����s����Y��sC��f�;�Q�qNn�:L�b�;���O*<��Eh<�ϗ�w��q�����;	���7�4��]����J����ƹWUU����Z�N�Z�xy���Ww��i�����I�i��Pj%}J�M�q�ӻ���n>�ܹ$\
7��kN3s��+)d��8��h���%v8+/������3h��"^�9L81�S��%x���?4���i+�H������Z���Q_O�$�R<Ps��b݇�>�a
�MԼ�u�/E2<���B��{��A���7�c,p`�+�㞎v�4G�Q8;�� z��!�[B�"m9=�_���	O���)p �q|����-�&w�@�Q�łn@�i#K�yO	�x6�$�q�]��p�G�!c�`p-�_���8���Y�YVPP���[u/{�i�G�jl���۷ڎm�E�9���o���<o���#����[�׋�̈ŋ�H���������?�~��_XnN� 0!�p�]ςݰ~�mܸ�W��Lx����O�T0�Q2B�u�m6h`��Tԓ	�k0�X|E�-��ow��~�z	��6a�*FÚ���g����Ͳ�s܃�P%��C���Z6d�`���sl�ԩb���v��w.(R�'�֩4 d�P�P7��;�C������0��:�B�CFȆ�����QR��BW��:X�I��Ki�!��q�lƌiR^K�(�
}��˩&��M<z�:� AX� SFҖ��m՛k��
k�Q���)���N�]Fz������Cm��aַO���H88.�I��V7�Gc����+O��=	E:�F`��2nڼ�W���;*ܧ8�32�}��x�1�M��<+�Shg�1���u���k4O.o���+���޹k��Z���6�P`8!�ɴ�* h�U?������PB����j��)�k��5{m�
c��Uh�Qt=�~5)(дPj[���KXJiAAؼi�m޼EJ�^�ŲCVv��?������촩�l��1#�8�2�E��NEDϡ�%B���1��{7.\Q�"����P8�*t��;�����<�����+�r��F��q½�I��(#�FڥR��И�˼�|���b����ãk�o^���;��`}+1F��l���N|��C����E!�oW����S�8�/mV#���0ߦ��\x�6z�h��2��!��(F�C�koC9Tq�$*^�q��+|�v��!��r=>��sY�/((��]�q�pxP�0����^�ݡ2B<�N�/� ���F�����Q�)cFI��"�>�զ�Ȃ�$7肜;f���'#v���]'%�J)���:&�
��:^q܍�(s�*Z�����  �I���b�r0���E����e��y�977��m��>G��SE3�0���Ϙ����������s3��B�5��&�2�YcS���p��#�G
Hd�x_�WA�&f,�?��{��~�2w�KƉ���8X���{y?c�q�X�)����A9�6x�F���O��V=��S4�����Z�yN������]�����v��Q;|�xn��Q�c6��A����ad�d;�u�u���/��Zr��0�q$E���o�HC/�L�F�p�/�0���4h�=A�z'pcH�|%���ʊϔ)Sܙ�N.q� �1�q\�T��2��d��F?+��9y��V���g�����2R�}�������$�;z�;�j�-�MS.[�t�J)��G?���{���{�LMD�/w,0�sm�k�N[�d�-]��(���-!M�?B��	
��A����|�.�@���475Z�6L�gٶ}��B���|J������7����%Y�m����{��>1�����ˑ#�m��U�n��[$�[-;O�sF��WU�q1~6�gfJ9j����:1�|���9v�ܹ2��
��S7��Z�uJD�8k���W�˯̷Õ�V%��#�*듭���R;���+��.��l���K-GF�T;���N���\�p������/[eu�e�YFJ���6�ߖ,�[T�'�Ij���-�w�~��w�y.�o���oڛk޴���(`�r�2ӯ_?�S-�(�(�̫�̴�౰Z��4)��+����'�0��0�q��W9$�}5P��C�66�Q͋c��m���ګ�K�>�p��T�Q�AI�(a��ꫯ�T���� G��Wd�~pRP^���c���G�	�{m2�dɨ�i_��,�7W-w��_F/�Uaa�+x�1���ϟ!5�F�(S���^`��f�/,-�WۢE��W^�;w��Z���p�(J
	
����D*��\�a���vy���v�u���sαV)���T�Y�W]�2���0�0v��~ᱴK�y��Un$�"�=��(O(]���B[x�'N��+��`VV�^&�r�tW�\v�S!1� ��G���m�6ON�$�$F�
Qh��;���P������VQ~��7bx��5Fs����U"�����z�|8�l���'e�C�pb� �/���˱.����۷Y���>}�8	��s���%7�Z�}ojzZ��D��_��v�oh�e���af/%�W��"�ǐ!C5��v��a)�u����þ}����\��<�����c�@���<q,�PU.��V{�U�{���8�����E0BRՏj�������^mu/o�p�[�.���K�*�rB�q��߿��ب��l��@���V_]�,����kE��vk$O�G@V�5o�ma<pt`����>Khg�]���m�8���&#��SR}�^q���}^P�)��H]}�UT�����@��T�PiiY�m!9U��g��ε�~�[��'>��m����7?�O����A�[��T3���/H� �ҿ������_���kTj�`��L����� ��$E9�! \v�ء{v�E�a�JyhOH�aÆ[�>E.$诼�=�n��f?a�����}2K�����23(��-�]( x�*���C�]0�.`�Q�[��^}�U�����+<m�4�ȼ����xF4�_���96���=$��4�+)j︉w��<*9�B`��T�����	KB%�T68S����͛6ٞ�l��}���֬[<1[J�+x�ۤ������#���k�ڔ3ϴ��[?	�)#(�A9��1O�BX%V.��j	�����XE��жn�a;w��W!e��-Ѫ[2��Y���Ϊ����%6zx��x�l;w�$�n[���]���؆�>��w/�opz\J�q)��6�8nܸ��vc5&�R%��dБ8#W�{0*+�ڹ�L��Cڞ=�\ �Cɦ�Q+ ���~�8�V�e�L�����g/�{�^[�n����:�y6^�z.�\CǍ�z���:�,�5k��2`��J��NHXm}�C�cC ���������G����JFB?JJƾ}��U�?����8H�.K�!(�̕����W����w;΀1�E#X\A�;�g��WOP䳎B( p�G��}��c�m�S��O<�1����8.�	��?
��/%�ꫯ��.���	
]����0��V�TY�#̌L��>Ƅ�I*F,���o��3��'ׁ	~L��̷��v_���6\s��v�΢�bKId%�B8�?�L��.�7흪o!��K����B��c���V��Q�r`��^�q�}��B������=�B1����Z+�-?/�y�	���}���̟����m-N��d$��cǉ��H�~��?�,�� 78`e�1%�O��i��� M�9˜nj��cG�\� *��s.�Ԧ�}��"V�3s��sV��NRN+�S��.�Ĥ,��e��m�a-|��͛7��DHI�O�9^&O>K2,��i
�w�c2A��n�륾�ʍ$�G�ݻw��@Zg�F����l�8q�J�>�v���9��}������h�+V�p|1?sƏ� �8K��y�9?��Y�9h�Oh�駟���z�q�����S��*..�0��.�#=":>)��췬=�!�v1��M�"��5�0�g	I-������������|P:T}ͷ���;���?�@
���/�3�����1�Q,����XA:�3���oE2:(;$���{�����E�V�8|'|c�L����Z;w�yv�g�9�#���~���s�<��!5=UJ�@���F	�����|(<O���^�-��b	r�t/�	!I,|jj�U�i��5�^��`�J
²�X�mݾŲ�3ݻ�P�����R��\e�!1��ʄ7�����;ڤ�u<D%#��aR;Ij����꿬���=~�M>�l۳��_�^J�h;s�$�8v�^{�9.{���Y���>�%�`պ��w!���~���T~�<�b�P>&%�����'��QL�-91M8L�&	Ai�6v�Lw��0E
Ui�<�:y���{��_[NV��Yc}��bP�!�>;b�!}u��E����((�(pu޷J���ԧ����,=%�{�Wb��Mv��^�{�\���w&��[����1
ȸ�B���/���Y4��c5* �@B�u㩥U8��0�|�h����QC=FiDE��
�aC�_��R��p9x𐌚=zW��s�0�W=L�a�n�xc��G�s�����R?0����2�C	��&�N4C۬`�R�p��8{1|��u�K[{�{����/&q��-[6�>�6IXia�BC�	\���#8u�>|�p6@����!�X]{L����Q�!8B�h���mㄩW�(�(R�]�D~�!�%��0� t�\�9�+{�'��	e�U4<��8a�D1j��G�V���L8����=��}�7��F��⼄�:��o����K�.��:���|	}�gI�<����P"94^xW0�B��E�^C�a+�=�P�}��[M]���M_��|ŀ ڧ�^*�3���o��f_4۾��_���̌�����\�~}4�%���s\99yz6������v�_��n*ㆱ�c��	FdNAQ�	�8=��K�O��(f~"O�����,�y�yv���[_;{���Ͳ�;�٦M���D���4u�96r�D��=n;v�v�~(�I����|a��Ə��ŋy�"c���쩭v\"9a�$_Ae�B��)�Pv�;}eL��
�K�J��|P��^����Da���o�
M\�t�ׄZ��g|X�d�r�Es����^�;�.�f�H��u/�\��_��,���W��g�#_��� \�ͅ�^zɝd����O��x�t��S�:N���{b;�Xx��a��Es-��<]�i�O����!��G}�V�Z��y�1�8��;󁽂o�'�5�yx-8#|<K� �1���vf����'�}ī��׿|�>��;�k��������O��@ZZ�)2��ӱ��-�M�D�x�������?���c��w������w�q����sVԧ�O^&{ksX!`�3�TLj�C�mR� ��/	J������QR^w��s��7�;��$a�1��
���{dN,e���X^61��
�ӢFf{##�c��O�� '%	�~��s��������_�}A�MMUMK���\1�&k�!��a�v��6��B��/x���o1EVZf�U�7YcK��7��M�l;��u��yS'�YgM�O��}
�{boJ��"\Q��@��p	��&U�� C�֐���V݋�ʪCZF^���a�rsl�3�l�1t�͘6�Ξ�m�G+l���#���Y��j���gcw��2���<o��-�O=l������w�W��qrJ��c��H�M�t���&��W_�	�د~}��3��F|�#�����dZFȀG�cA9�aO��:]#��
fpX̺Ka�-ى�P�7ـ��k��}>�=�����]��&aK�_��q`tq�}V᷈�x-��au����|>�����<W|��G�p��s�E|���B���*������|�]}�����ו�~�X�g�N_�wx`IV NP���Ɣ��1��y3^�h�w�WǙ�οY�c�i����`Ɖ��6�[��P���B?(����0(S�'x�Q �R��	F0��g�C"c�����A��\�}�(��+���`\���Ǔ��3f8/�p��'�7m�����I��V�é��ɢ�I^��A�I��D��f��W��>�����/|��S�_w�9|О~�Y۸a��;��#�_�ڀ.x'G;44�줔�/ǳ>O�[`IVX\h3Ο���D>t���;���mTY�I7l�]�v���-O󸿔���$�+����r�f�!a�ӧO�믿�V�Xi��w>`�O��P�xR�eŗq�7��@r�*$v��쳩�m8!w1*Ie30�t~h���+b������&�{�ej�{�����Yq� �<��������+$�0��+�}��7θh��_�)Q}#�Pp.B���=A8�HDaG��������~-ڥ�8�<��Dϗ�ie#F�&�8�O��������b���a Y@��,d��zr����K4��N�-�}C���3��OBjy����B����M�*op@5_!�#��;�M���ϴ|�v͓Eڹ��_�A�G$�+��կ~������&�[N�����6E�t�ҥK$����R.'�o���I�R9�ҳO?m�8Å���b�OlB�`V0� LF�ڞ�=EE�Y�_xȾ�o��|��u�������?|����>E���Mj��2L���0����D!���a@T���Cq���F�!�G�>��ɧ���]u�e��/}�~~���N���;��%4�bf�x�`�l ��&CIx;0w�^9Y�s�{��/��a��ĩ2�*�j����a��E���=Q¡��8��U������.�k���G�%ˬ�R+��׽d�B�	�-�H�)a/l4���nJ�����S[s�l��)?1�j��^*��Ȇj��)v�.ۆlgNk���#���϶{>�Q{쑇�W�����F+,*tFO(B���+�W��ǚ��~��R<<�p���&��W�&W+�e'gZi�ȹ�^�|�}��O����&eæ��=5�)?;�L^/Uo�)e�?*+�4��(�xQ�|E��V���5H07Yzv�]6�R#$���|�3�&� J���Q�.��r��o�[�	e#&a���G�G���&�0���� ��<>_4�u�{`��=�|n��F�����_Ƌ�LEp�l@�ذa������>�*�Cȵ�3������8��2�ߧ8E��L_�<�6�}���PXMKOO�2t�C-�J������x�I��=A��0f�Gf��A�<C��>���'7����|��x���D�)���+��N��+��������FOx�r���,%H��=(���B�^C�ӗk�[��퓬����
�1����rA�>���^Hj�Ӿ��������X������-�{R�7,�H@:L�Y�a�У�c����k"���#�K/��x.�ל����ǎZIQ�mܴ���_�x{�-�2�d�"�g������$�`����ýǫ�{��{���b=�|�}荱kn�3Θl�%�&M�`;�oל����]2P��Ъ��i�����3�E��waP��/�0_�U0n��s�o�>�"NH$�d+�7p�ׯ�h�7o��ڲ7�9�QR|.�9^�Ư�Z��!xLx�;�3����>)|�KV�ǌ����!��<q��+�O>��=��Sn���`�2�.�9ӏۀ�@G�8Vf6K����!o����޶hL0���\V<��0���1�1"�k�O0�����ϣG��������	�C�'�Y�=5�c����:�����Ѯ�{��Ȳ��>���֊o���|�c��t� �{�i_�H��Ӧ���/e�׭[7��7��_���R����G��>����?n�ǎuF���bCw�>S�����v����[��SK���+V�f	����_�׿�5��g�A��g>k?��X*�Q��#]���'����F���Yا��B��-*X�C���fVV�n7�x�Id�[�l�+��/,�g��ͽN�o��E�����s�J�/�'��1kj�r�Mh�|8� 	�XfZ�ÏW�Tw��^d��I�m��v��ڎ��m������ex�Yf{�T��K�^n?��O�B����-Z�����-����B���>cØp>!?0a
p�rOdެܱ)8+3[Ɣٱ�jKHͰ26L�X�����y�Vߛ-?;��R�m���_`���ږM��G��۳�ͩ;D5�\W$H��D(�Dw�P�_�G�(�^B��SҤlNpF�DrJ��1y��;���Ά����xR������5��gͶ]Rn>����3O=�c(n����Ԥ4)A!�BG���������n���V�z�}z�5UV6|�ͽ�
�um�W�|�KVc"�ث��G�{�TY��}��~v�СC�S����X5�,������.��Q!xQ@y��;��s�r��y� �=�B{���'�pAΜAQ�X�,���g���y��o�(G�0F\qmaxQ��ڗB+}�1f,�66���V7(�,��2�8f��q֬�x��~��m��is#��r�c-���.:����+m�aW���/�W��u�{�1�y�q?xF�LI�:� k�>%ži��A?S-5َU�I�3��&�Y�ٱ_��W�{b���iz��%����>r�.���9�d;d��h��ø�h0.�����/>��y�{�1b�}�B�d�o)�3q���O��@f8BZ�oV�3ںm�Uʠ�8Za�ϟn���o|/�|������C=��/�I�,Y�K�@���;�=�U�#��]��ap�p�{�CT�,vC4Ǯ��*wZ����*DZ�L��;���Znv�=��ö[��P�,MRYC��G�%��L��V�JM�h����x'� �@��!��{��^{׻��0�O���Ga"�D�S�g����!X���s��l�<P"��<�0�����G)�z{���B�h�O�"�:eUrD�0�X�ȋٳg�{c�<^e8\���^�xһ����
ש��P`�%��,�?�D�9�p�x�w�aseq�|�T��R,��=Fɼy�lɒ%�_�r��*�
�B�����m )��qL.`�;�����x�S�)8�;���Dy=g��Ky���I���$�՜'��i]���᯴�n�z��O�����+oT��_=h��Ö��q�����������[N�$Oo9mʇ>���2f����*a�/��������'�w���>��,s��@40�����t�w��ac��}4�ɦ��UH�=f�]~�庿ޞ�9	�"1�Kt�^O��%D� ���&A6=��4
� 5�1�_�	�0?�-鋧L���`F�?">%��y�w�����%vδsmݺ-�n�fKM��'����2���=<K���@��
�Dx�>���*�*�X�Q+=�n��K����52�Ġӳe@IY��
���<N�[o��ŋ��v�J���|��ÀĻ�P*B�������aea��@B�TV�Z���fY٘q�-M��ۘb�5G{��Sf}��lT�kmn��G�YC��K{���R��y����������#
E�d�CŘ�x�a`?���w��!r�eWH	m��(�W��SRDKJ
��8_F��<Ѥ�gؠ�A����˾ј.����jFGP`��s�c�;c����.(���v����ӟ��5�������Ν��^B.�/��ezG��������}�s�w�Ȅ���.�S�D$ |QT�<����jܓ�a���I|s�ֶ63�aa+쉙8�t�ɾ/�e��Pr�E/+��o���%���#�0V��g܂Ҟku�a_�����{��'i.	�V�ι��8�Y�.�����/5��7�g������ɜ&�x��$���G��c�	�n��oR��G��qp��Hp�����Rׂ��U¬�J�[�n��}���-�01�ehV GV"����0�8/B�g�@��mO̐�X�vp����x�9��a��df۰a�Æ�
-3~���EP�ڂ���O��pN���e"q�{�z���̜5��>c�9 ���w����0���s���f��	E{�~l�f�0��cE��W�p��{p��=�~x	��ݯ�=�<��g�}�}�#q��ϡ�ր�1��[��nt<�*�!,x5���Ul֕�AD� V�5p>?�fQl��>����#�K(|8���Q�3���1XP��t�1jB�'�Ca⤉v��|�x�̎����V��?�5DU@7!l5�|q�8�]f�1�#G���s��8ײe(aHr^�@� 7���c!�<iϑ��W�%�1t��Bh�^"�`�]�7��@����|;}dlY����-��|5>��⭿�կ|ܙg�)��Y�<�C���{ƥC�t�Q���Uͻ�@n(��p�V�9|F�G+��R�����Q�Fۭ��j�\r�]8�B��۶n�!NJ��g|�od<I^��G����_me#�
�d[��M��ԓ��T#Zz�쳧l��׾����w@�5�N�"��"�h�����E���+����
���x6o�j�e���(�4�	wA��k���vۻ�hz��<�
*6���UW͵+������?��i���6b�-�R��x|�{��lI���T�?�9g��:��apݙb����^�#F�,1�?�d7�1z�I�K��۷ZBj��x���K�-c�~�U�x��v���0P��LuA���H�r������b��#�DC�n��������EK�x�DRJ���Y=��xm�q��+�?�Z���]7Y���W_y]8j��@�)S�JHU��}�W(z(3�F��#(0rE�F)5v�F��%W\i�%t�m�l6n��L6�g/����,��Rd(55U[B�O��U�o�d�x�: %�?�)�����E�G(ˌ5��N��xcU�����$��o��n{�{m��7l����V��q�����Kv������y�&W�Pl�>�iaF�{H����c�UpA[���x٘OA�с��+������[�j�b��"B��8tp��N��n	���`.��'�<���RNn����(��3��s�9l^4��r��`�����D$�h#��,�_P�Ih���cƌ�=��ʕ+��	t+Z�6x7��ڵ�ԇlKİdU(�{0l���	��~Ǹ'�:+\G�"�<O��/�+�2V�L_��޵^��P�3�)�.)�w�����T}1�&xG�w�Y��Fyw#'��4o�Y�醒>�RQF�Jp��I;�gY�,���|�PpP|���
)��{x"��9�E��qL����[�d,����E
ף��h�J\F���|w`�8�;�R����'�Xc�:(|m�b���(�x�Qj/�4������
>p�w*)Vl��Q\�'�̞}�;qX]�z������������8C��Y�b�hs��r�-�w�~[��j�1�y7�;{Ax8NEα�`�'��0@��s�(��>Q>����m����z�a7"�+
.������^P�'8 %ًƪ	+�ƧC�<�H���M%�q:�'��5���m`�ޘ򙒣Dn�/�]�+n8ĐO�Ŋ���=l�Pʊ�
c����r"0��^p��]�7�=�76�:�����d�N�>æ�{��G?w��Ȅg�>4F$�!0�8o�$�!x��HS��������G��sU�
,������#�vδi6뢋\W!C!	��d���.e����>���x��fO�.��@b�l��d�S�'� vdw����!�	���Hc�X�O�6�Ymd!�:�q�s�0�R�>$�Ag���{�.�G�-̽�1�ࡾ������D�iv�sm����]�-[�y�)��\}��?#]`�#���#J�����#A�=M�]O`JC6���1q1�Zkjl�)�N�9��!�a�0���/��ÿ�0w�51�������gM�Bt�������V�o�[q�$�q�%z�̚[S��A.�$b��������2�g�0X�;J���������"�i�z1����W�{7���`!P�>b�\�Y���j��ٔiS-]B��[k;���@)��o!���ٹ_EpR�@��B�%p�������dC�N�F���4Q��˭��Zl����2 몫l��mf����sO��={�9RBf�gy��5��E2Bkշ�l�Ν.�0��O�W��G�����P`U!]��������6ML�C�=���~�r;�w�mX��mݼ�d(���۶J��)%g���2�䍕���{�n1nV�6z���r�PƆc�]	�'���O�ϕ@���%t�dD6��L��o���]%#{����k�:۩��R/�J�P[����;?r��:ڕ�_������n�"ʌ9�I�U-��G�Dhz�`�x}Y�C8#J�+	dK�>%E�����/�c�=���m�WI��ہ���0����~֑^�Y9kj��P$=}����f{V�A{_z����A]!-{��y��A���j���zH�DZ�%k\�2��Qӻ#)�c���b�J[�r���|���w��i%=5g��&�{�YeU��^��{�a�)�GI� Ƹ)MxCX'�q��
�Օ�������{	y	+�i��9��qJ�ȱ¾�lȨ27<wlߥ�Hƻ4�"8J���޷���}�<L��x�BƜ��a���'Ƹ&�02;�>9�EJ� �6)��j7C�f�eHՐ�#%��3}�yR�s��p pH��3i�<�,���l�UWX٨��O��ص�~�����7�x�O�B��b���V/ٛ$�D�R�T��^����臌���!�=B»`ĸ�ߑN�ߡWV�	Ձ'vG�?>��O=��=-����pl��������0ꙇ���O˕G�0H"�T�'ExB�%�s��0b�|��K/�UtR��8�<&�A�qfz�͞5ۆjSϞb_4�rś�����`.}�K+�=��+��#'W�4:F㏹�,�~0:�/���~>�9N0���q���Зe q�u?)���h��Cŏ�;�6���C�?�E
7B��fff�;�С�Q�֤��Z�Ǝ�g$����%���4�fL��E�'��ì�1����B�Ɏ�q>����8d<9(�bh�'�����?
c�5x	�rF�n�dZ��d������g��3'ۺukd\�)�2Ԥ�'�Ӻ�넣z�|�v��pɫ�R�_{}��V�g�#|�D~Q�eJ�Tw�����'+���bA������+��28m��)g��
IJd�-Y�������?���#�Q���o8q�0��� 1�=��{�}<�-�T���	h>:_$~W�O&B Xhc�}�ی�4�:m����1�n����2�6��Y��}���I�y��ÏH����w:��� 3�p&&&�Ɉ
¶��c
<���&E��533�M��#0�&�� ��9�b��}{�X6{��`�pO)g#�ܹ�3#�����������/t��&�1!�0���'z����ߞx|�=��<��>m�R6�3�o��_Xj9�},[̫�-&�
DJ��M��#)͢��$1.	~���(�|!az������������W��[ԟ\4p�]yŕv����ޞ�a����ʳ��G�$Y?	ȴ�\1O#^E���q��u.��V�Pa�k.��&&��)<"�tE3G
�P	4��5����l��3,[�mqn��[dǌ�gL�ϟ!au�}����|�п��K�ӯ���9JIb�x����+��d�E��pRWp��>R襨��6J�>��D��c�S?P��~�[[�꫖*!5z� 8�C��H�UUTY��c���l�&M�s���sC,3?�ʫK�>�q��E�A�� `e@mu���`'N?Q���~7X�ҽ)�YNA�%�%X�OF{���F��K��-α�3���ŅYRۭ��V	���O�AA�C0UW׸��[�O1�_t��hX\���ce�ſ��ve�Qx%d-�q���(E��瞵������.�u���]�p�+c�2Β��l�������JX/�����1)����Cɪ�j��ZVs2-G4��]�T%H���Ek	�R<�ݰMNK��-e��J���Jy���*��Oi��s��6H�Kq�>6�1�~���}��r$�@�Cq=v�/)�^�{`FJ�6|��d/s����~�U���u����a��O�
�ꎕ�\�ڜ(�mOL�c�uV'�&f�ڡ�G�J��א�疍�����"rÍ��M7�䎗7�X�mV�x7+e��b���7J4�vhKd冓�HV�ɰnwE)Y���ʰ\͗cCm����˯�q�&�ƍ��@�N�d�E���zz�S5�5ٙ�x�)=��sϱIg�����
~XI�����$>7�ߪB��O�Y*ʡ�gvF��9]$t���B縩3ΒÃ~�H8Ç"�@S��Zc%'�5�L(n����Cj�/`b^
�z?�Y}eK�Ą���.�C�xy��
�'e��a6��'}n��	��( �`޼'��>��/�Q�&M�1��~&�vx��}�,�)�Iw.8$����_��v���EQf%~C��7�&�'U$�9*:��`�ʝ�I����9�'#�o�n[#wㆍn$��!�q����sA�!v�K4�����;�A�֡���u�X�Rݙgʛ|�d_M礵9>K���H�Vڿ�J�NL�pG
����ύ7؋/�(:{ͣ�/�a9jT�� �Lj����/*Q'��KS�%$�}xm2n����F-�agJ&��i���O�C4v�{��t�L�A�Jݐ7a����+��<yR�tޝ��/c�Dr=�WqY}�-�q�o
�;8?�-��8'XmceÆ�٧��;i�D?̗�I>2�_?۶u���W���K�����+V���ߨ�vVe�]FC��M�U�o9��_b���"-5S�%YU%GT{H��i�|^a��5�ـ��܀g��5��0���k���/m��ź�mذN��9�d�d�+�ZcK��+��98^�p~{�|�DӬ��SP�Vt�,X ����
���&�_�Z��?���DJF{�:�L���rC�������sˤ���3������6����Ϲ�����@i!<��_��!62�@������ٞݜ��!Q"F����a:�}�q���T��C�x�${سPV6BL�Y0��Q�[�y 	c�OB��Vt��[�j�=���f�KE��{��k���r��i����"0�gX��]Q���E����R�߮]{m���2X�}=�<5��r��;>�~{׻n�������f�װ�.�O3-U}��'�������/6�3fx����Yԇ��I>��c����Ϯ��F1�=D�{DL��rx�7إ�^b'���d��=�2%$��.�HLzn^�{Q�HŎ�Ǳc��MĠ�z)�U	��h����Z���?�����_���a��9<�Rv�����r���#G=�	�l�a����T�]�#h�q�^��ac��t�wE���ڭ۶؈�e6s��v�5W�̙��\��Ɵ�����OoeU���ҋ�ꫯٺu���V}�X�P�ӨN#��M%r�3V	�e�ȑ��*�-�@
���)+�h�;զM�l7�r�͚y�{>��q�O�@�3����w�J����=v��w��c޼�l�f�����a/-� J��'�W�9�0[
��g#�43+���{w�x�]l%R�	�B�a~��&�p��ʗ��y����?����'?sE�d��/%�a����g�7n{IƔ�D��-<�G���>���aE�=�x��S���D;6l���=��ph��cՆ�[k׭�-[���(x�;Nį��9m�P����9/&̋#2�<8�>V����z�|��x�"��=������f��ɞ�8� ���� W�@B'���;㧺�96����B���m���b���Kp���d�awl�'l����Ͻ`�_�.��+�:d���BƊ4��O!c���  c�b0��������B�p���n������r����@OQ��M��K���"L����0d����-�p6��(քa�7���F ���cR��7
:�ٛ�x��֨�
�r���0e��_r~�.�����6�R�a�(�̷sΙn�D/����u���0:�m��2F(g�;
�>b����M����w�i�S�a|"��\��
Q��B	��o�ɽ� O����������cFX�_<���8����9d'���`�y��IV̐5�վ�x��{�p2�g�d�x��'ƞ�q�+Q.�m���c~|B{�G���v����ɰn����Sm������U����̙��#�<���-��k �f�ӟ�g��ݻ/�@)��2�a�0
����P*Ia�;�I�ۿ�[���k��bH�E>l�3�|	�p�K�3ob�aF$F�i�{r����ߊil���V;^Qc-M�Tq2�55ֻ�e���fdV�F���&�;`�ΌUa�O>����o����/Z�JhО=�e0mw��uk�����O�K��j6�F)�(t�Y���d	�!�fƻy_�"L׉�'_�t'x�	�IU?k%���?����˃�[��.\���c{vn�5k�����7��+/�bO�{������駞W{�o������h&'L�1��IE���-6��7`��j����	��T�f_}�5�)�x�
Ye�͕�e�4IH��̇����=���2<�����d��lڸ�7A���wû�J���cn �նX�w��C��'������T�Ҹ�����ߴ�o��7�Xa-��;���b�m�f<��c�ʀqD���_�����UDh����G��S	�����y����w�NI��w�?��v����;��`S�N����r�җ�l���Н(0(��O1Nd	C�Pu�N�̠L�:�ʪ��Z��SO�gZS+��e�ej�jl��]�{�v)[{m���k�ۑ���-l�F����t�<��D�?���+��0n!˕x�H+�͓��
s������cG���K�xx�૭��Xkɩ	6jt�M7��%���d��^t�E�!~}�k�����(�%�L^n����h, �n*��n�nVΡg�DV�8�lD�]w�u�������W���� NF,x#4��5^�t��"9����f7�QvP��U��2?G�R��� j����9ٙ���j��*��F�8�h�;$��X	^'㌽)(��O��%K핗_�߁�ʘ]s�5�`b������(�3�������_ҧد�O�@�D��1�>��^���ܹW��>�9�E��	c��(�rƆ�Q�;���9��1�'8����*������L��PZ��3�;=�Ghx����
6�q��*�0c�o�MpW�)�qsR�X�z�\�J��"*yE���&:\(��}/0�ld��^B<Ǎ�:�ߵl�~��=?(��8���������w���g\��[X�i/�O�k�(�x�]�� ������bࠁN��͘ ��\@W�ė_x��	0£
.�����J�o� �'mE�J4��;�X��&����/�{i\�G�:���yW��qeL1Nx�灇O�)X��:}�_&���*2��
N�%��s�4�|�d�	��}g�+e\���N�e_�~8UH:�XB`��3���<�+�t��hVV��t�u6�t��O��~Þ~�)� �R���?����_�zo��wJ�5�N�r�=w#�LL�a�W��K/u�C���f��(	0�q��x
W
+L�G{̙
�v�<u/�L!��j���p�"o���W2J�Y}m�ef��/܋'�$x(10<�S��Yu�0S*���0H)Lc���!U4�~)lG#��|�]�� �BJ�v۩���k%R�ɢ�(��bQB��*�Y�,0��խ������#!0�Z��o�Dz��E(�P���Ƃ2y��~1�r��2a�X��{W._*�xH
S�����������hb$q`*�	6|���1�-x��L� ��''[�K�̑�R�,�_��W��c<�m��Pd����H?���mi��X�آ�ʠZe�U�v��Qg�d�+9³3�oڴ������'8��� i�}bI�[��O/�˖1}���v�~��Ql���|��.��|s�]z�ł��=ƻw�1�q�hI�~nD#����1b�z�8�Q�F�a� �XE"4�P���2�ް'd���@�{�4�}�Wƈ��@�^�x��
-�禮�^oY�8�C���]P�(1�B(gBB�N�,�t��$�Y���p����^��y��X��K�N���{Ą�����O�3���^�����K���Dc)
�q:
s�1������Ϯ-c�����9��Ԩ�dE�_�O��֬yӞyb��۹k�?�����r�J�E��?�~g������-�W���1�Q��#�}����߀�1F8���M���/�w2�^t�+�(��#}�păC�M��f�^����~ ���h�����,�ԗ������i���|Y��aU:��?�0�͛7��� S)`��(�#	���f)��d�a�>��'>�	�����8���\QY���m�$�$0*���<*��!�������<��p2s�L?��~�����CS�G�s���I�����d��g#<���K��D祌;��g���?���F��:�J��h�����~�����n�!{Əq#���E�G�%U�ɳa<��~bt�;d���� c:e��2
���Q���N����	݄6��U|q�0X)��t@�2�Ƚ����e�ĿW�\�����9�@��f��(�x��� V<����:�,������s�w�3H�ĘaP��~{����g�q� ��~㘂K�!tL������3;ڀ_O�:�i	��cJ[�4P�8����~�z76ῌ��6��\!L�3��"N��@_A�`50G�{�vι�����8���p��J�S�eL�%Nx<�p�8a�D� vj�Ɖ�%#+<j��y7��_*\��f��7_o�@J�\��~RS��f͚9��3������K���Ӻ�H�Y���>;LJȥ�}c���ɉA�QV�0�`f�a��&��C9S!��G�h���\�J

����@Ɩ;������_����cr��!Y6��%(3��֒�K
8Jrmm��'�NP�)Q(ſa���!pal\�=��_���A�vᬋ|
�
�>�j6c�yR�rm��7�������7`��1�LOb �8����*����y7�w���y$�/���5d�`7����a:���:W:��3�:)�R4.�l�:�C��5�m��֧���"W~��� ,��C����W�`G���r�itiVSW�xG�ƴ$�*�x�N�  DY���?r�h�R�xz(E�0�#��w��	z�@���;H*ѯ_���\g{Hd��؀~�A��x�P�X�#�[��
a#l��X�) !�{zZ��@��E�����W2��ō@<���Т�W]�ix�<EV�����c���>����P���"[� �%×�A�ęG�B�e\���c���M���^x
�wVu��
�[���d76����~�#���~Ŧ�3�V�-�3^a��Aa��ď�v0Bsdp�=%$���*���U6&�1�%@�w���_�49�F?���S�F�zW_s\��d#�FH(�*q�
<�h����;?�1#ԛR��Z;|n�����k�ϩ��;B���P8��O����/�q�����v��o��ϒbq�{JI}�e�����m��2�'�.�R���ڃ�� �������);C�a<p|@[�Y24���+�g,(���~��@H&��ܵ�U�:BSY�?�� }d������P��K�/�"�c|0��A�U�#r���d���$&W5���B�Jd_�}M��pH�%
���0����Yg����6B����{0H��Y;q���P�p\<#z��|�h��(�|ҿs�D)ɑ�ʴ�7(��&��/��F�s�vY�|��G�\��������B�K�p��|)*ь)0D\`  /�/����;mD�wVm�.��1�i����1n�3!v��h�B�����yƔ~0(���@���V%����YV��{3�Q$/"s0���!	�0��t�Z2��~Rk�78���	|H�����%Ii~��;��}���'�@0�)$���a�����*(xc������AF�ߟ~�iKVk�#8�i����Cd�1((��<�c��W�
��;c�{��.��'x4�~��h Q���lD����ٽ��:�D�x�n�F�"��� ��<�A���'N[�(��������ʠ��}��e��� @���f\1����t�����	2>��E8-8���@�x�#����km��z^���նh�Ɇ���/����g��V�[=~��,��iV�3��ȑ#}�|�Ζ}�;��~���=5&َ�Ν�'g�S��PI���K��s]x�{�,Z�E�x���ʫ����  �oIDAT�O>a�֮��(f_t�X��J�f/{U>("�V��>UU]��	�oJdЄ���`Px��h�����d�G��Ig�iC�wŋ�`<�׬߰�C��$��3��%C�
�RFQ���T��pvL��)|��77c �����C��i�f)t(�x-�������ӟ��B�g�	!\��� ��o�۷w���s����AR�d�H�$W{����a�*�%+5d��]�QP��@J��3�F�� ^�9^�iS�yV�6Ayyپb��V,�`�!8�\�R���<3	�KH�^���K�@��$��`��˒@,�1Ө�׸��:ډî�+V�B�FD=��s�c�v$�^~��SB�Z�I������e��ݐ%�%
y�g6pR�qB`�d����t�/AJF�Q���JE�a�x�:i]�	���j֍XA��]a6��ݬV	S�N�3�H�@l��m�ሲ��{��Q�olv���C|N:�[�V���c�k��ܬ<�l�ǘ�` 0/9H�b)�̧g�^4�dÇ�p��
�<�|�o:g�!OeN���"�կ~U�֛2������ε�_l;v�]��:~'�K^(e��?�A_y�'q�-!`(��N?W�.��l�C�#��Kf&����������B�'��;��h����ݗdÇ����W��+�
J
F$�߆�0�.��r�Z���5k�ܫ�B�BJlظ�V���� �,�N� 3|�UV����S�~�J�!�NfUנC����w2½��w;'�6پ0�P�c�$G1�ݳ�ߏ��
 +P8���O�{��GgFeg�$0Gc��ADp���7NV��uB��<�瘋�� ��Eqd�Y|���?���>���G�Y>�i�.�߂7�|����¡�(����|�b�1N�V��8x�&�����J�q&���U����0����&���*x*a�D;�9���<�8|9Ī8��jC�r�����i��!�w�n��G���}*��a0 /�A�࿓
F9x�_3�1x1^��1cE�Ӆ�"7��>�u�~�z�-��>N�90f���?���n7���k�6�=ࠂ�V[���X@Wq<Y��@�L��p?�W�7h�+�ɼd��q�}�a���¹���^w���z�o��+s��I�y?4]0�(a���D��&*+�-½l�R�	�M�/0S�g��9��}��9_�(*
��a�s�!��R8�ju�"#O����\��D��?;;;�n��:HÄ�d�ɻ�4o�kgϞ���)SW~�k_�]Az��^�4+w���2)Os�d�@��a�tP`��` ���K_��3R'#zLj��xn��(�+�/�}��f*
�<$0/&=��9�H�u��.x0��XD�˂�<;^qL��~�B*Y�*0A��1`@���O���4���!�2�9�1����l&fS|mu���\kmjs�n-����vP��/�6x� 60w#}��Ge��!F�+��b�y����-Y�mG{�q�567��R������:�e�}��}���,O��P'�_��{�Ȱ��W f�i{�<����{��!�#+�O�/�K�C��^XɁ�7<���}s9�HW�ޤl���{\��%�ђ���_��;�zo�q	�M�\t�!��{�����A�����̸"���5�υNg�F��Kx�Zy�Z��F��� �QSU)�C�	w}d���+8�U |kVe�ZE��>�!�8��r.�1����P�����R���dqIzz�������M�6�a`%���G���.#�MW��;���pE��*��<������2���<�aO��"Z��	g�p�c{� w@����>���wYA~�͘q��3�LLu���9�"H�B�=\ol��>^'a�+��\�B�~hك~��>�G��G��k��/>Z�㝭�4��d�a��N���
n���@�A�g>��� ���ضu������d���R��[�%?���$�qg��-�&�$�p�F���~�J#|��\�M;���a>�3?������GM�Vx�m���/��{�Q�����B�R��IxF�G$h`��	��HyN
x`�����x� �4a����q�0%#�*�Dᅷ�ڵ����?a��,v���1"� ��Ç{�sx:�R�y�^��1�~�կT7"Q��?ㄳ�U4�T�UƓ 
	��`���a ~��a���	�a@��O�M�_�No|B[��L�~�/c�.V�H��81���Ϣ@��}%\vy��ˁ���o�ý��jaS?��p����uPۿ|�_��뮵�^}�*�s�u�����TZ�|�s�W<X%��t����'h��8#�[�/p�F���aÞ�1���>�-�5;���%#�0�R��Y��s�5��X]������F%F��N�W�d���/%��X02~��a5�OV̐�q����Oǣ_���!L�����څ&�7�w�g�M�q�v�m9��ӟ�ǝ?7�t�]|�l���ř�X���]ډ�:\!v��VV�	�v�Gr�U�z�D;��9�� '���}��%��<�L�� �AX)�g�w�,OmBGT
����q��ڭ��h���5�G}�'��C^xт)S��ٻ���)��iV>��O���͑�RB�<�
 ��>kV��pε!����/2ձτ8�g�{�ʏ���v�Z���I�S@i
?K\iDx_=�
��'>f�]z�]z�%6����[n��瞣v�}�e��.H��;�0�VT0`�03<e0�A�9��%��{������e��M�6��+Uf�i��_�$m��ٵϦ�9پ��/�4)��z�~){pE�e�`�Df��
��y�}��B���lNs�s������`?��I`���[�~��xIQ!td鲥R�iT��#C�()j#e\nڸ���2ȅ\<������ł�cOCIIW1j��tFӾ��;�Ԭ�>rPp��@�/������ k�I�\C�8�I�H�p��k��B���c��`PF!+cX$��"H��K���s�LI9SWd8`T�7Lc�`�[Y"Ń�M�M�@�9BΪ����qL��Q#G�"�1Z�>l�`W80L��QPS�w`�����0`��d���+/���}aMx}-^�`�X�Ž��c�(�(?(Q8���p��烑��Ԓ�.�{g�J���p�dae����2�R��J���D8O�N�C�Z����fL����/����lْ�2TQ�����SI=�y��V�Yc�>�lg�j��~N(@��x��V�	E�Î:���D����(3��aCGj|�m��͞�m�Z���7�ҝ��Ij��y�f�m�@���]�F
s&�AB���Y�;�JҸ��	ZC�g�B�N��i)��2�2�j
����";o�y6f�W�Q�0��(�()?��O��Y�b���	{w6���* �S��E
uPAp��XAON_���(`"@w��R�r�5C��jj
�m�#RS�B�C �.�"�
����G�B���ڽ�sY6�[x'�yB�Q��R� |�;߱�|���_��۶l�(b-n�M9�,o��o،?N0V�Ȃ��2�}*۷o���<?�أ��K��F�O<GbpE$+���C�����$��R�#���w0v�FAp�����]� �R�)�q �B�K��������n0�'OE�6x?�9 \�I*��D�_�頻W̹ҝI�-���'�3R=�N�jQ�_�����@?|��iRK��`O0{���W_u���W^}ŝ}�Ř�ՌZ���H�@w�
��rġ�!�D��8�X]�hz�w�_�
ϳJD��yi~ÆM~@2�܎IF��c�y�cbp�+`��\��JH<�0>����Oۋ/��}�70��2�����x�3V��'��w��g�y��އ��F�8Ɯ�����	��;�'m2GqF!?s�k������5�X�*� ��I����I�*�֭]o�;�C��XD�.L��P2C�w/���fꉞ蓯vouM������~w�U�����K�K��5��9��@:���w�=\n��ÇJX*f�3���d�>��#.�'M+f�&&���R9�J�:.&�l;w�x���s�y�ː�%x��ܽ{��]�aLt���#l��& ����%by�	��[�n�^n^t�]6g�������0?[L<O���3q�|��Gj*kL���$D���U 7���_zQ
�)���kmJ���k��[^~���N�����9�\W��X��ʏu�j�����t}_��W,%J����@I�2lq�쐡�<='�c�=�+4(���7}�葖(k �2�o/�vdξ�n��f{�_��.�p����wҤ�,����\x��GP��k����$��ÙR���}����?jw��Q�s�l�+g\q���kj+��:�������ѣ|����ڀ�������y�3g�]~��6��i���K��������ʻ���l�5x�@��h�+*m���{�%�0xQ����'� 1b�>̶n��q�(�i)�_�pA<��*(�cƎ����vϘ->X4?�CQ�Hn��ʔ#K�����e��NXc��8G�\4�f}���������E.���($زe�mټ��XA�£�7eg��6NFp�=V���ޑ/�b�g�#� ��'|�����j��Rj�����0P�|�h���k���>��٤	�|2~�Ɠp�-[7�Z���o�G<�'M���@ƛ�
fr�+L��/�̳B�<Ŭڠpx�g���5p��2��m�����]뫩8L>~�v��W� ��͞m2.HiQiE)�{�W�%//x`����g��o������a�����w��傏�<�$�h��e�k>��h(��7���w�эک����!B�P�pT@��}���O|�㾪D��`D���6m�͑�@��2P��
_��KE'݇q�I�1��6�sFcN�{n�սރ��,�p�%Γ&L%ܴZ|>�Wc�yM�{�8����F���!Q {��`>Hs��o����%E������<C���ݳ��=�|�}����ÿ1�X5b��1��x�R��k�n�J�H�A_	<$�	���k��\$��F� ~u��9r��h1*ѱ�;+n�n<�Fr1,ۅg�8K�mi�qc&��ٽw�;N�����-dan���C�G��>ƟU�/(�m��I7�GU�LB&�+��j)�Wν�}5j���E�΋�M�2l&��gM���A��M+����z����@��كܪ�$�y�M��k��&����VbR�����O<m�_;pp��t�m�Y��}ј���S�B*�<�3x�h+E�7���<���#�3yb�'�z��@Fέ۶���2�22�O��`�klCx&�� [0�w7��KY���96k�L�g#N�#G��^B�S�Fݙ�O�&�6���e8�p~�o����1OT��1���BȻ1n(��8�+\q���pg�ޙ��y�VRT���Q����#���p�>�裶F��(�q��< z�#�)��}��;H8�0�q��[b��z���)lɶf�F��w�>j/����2�W}��i�{�i_z�Ӭ|�3�v���K������&��؉Qq�Y������Wl�-�m����{R�� �d, ؖ��B(~���w�~�����wJv%V4P��x��0j�x�~C���:t��ܽ�^������آ�mذ�Q�c��{s�a/
u��BH�bJ�FJ\1VdS����F�c�)�c�x���d$6���;�j�}U$55Q��oi��|�'YB�sH�v�D�VL0���Kܨg$fH��kþ�!CJq)p��]_�2��'����S��^��p��.;����"#�M�4<�-R�R_Ιj�G����t۴a��.��J��Q!AƘD���$EA�F�y�E��de����J��>��;]�#�/�eK�T�"��z���
���{��m�q�F�����������y��x>b��D?`u�fHYZ$��.e��E�(����<
���ˌt���ӄr���h�y�,�\������G�!rH�G�L��W���n�=��<)��6e�Y2���ꫯ����ӂ�_�ўy�Y�%6Ⱥ ,T�c	G�oj��<;^Y.��!�\8�������?t�Ʋe~F43�t�+�&qB��/�,�w��(����_;���^�B"Ã}#��0�Pd1k4/1��� ��"��T*ս��ϗ�x�=���&����TkK�,�p�;��<��M��8����A�0�h <�Jh��2`�,\Μ5�W�؛n����]� �M��/��J���<)��dq緿�M��]�ڠ�~�l�B{����E���r�҅�N8#l옐���U�<f#�e�}�]v�m7�豣<%��mƐ61tQ� N�����F��Q�@#���_��]>w�;/p��@X+\|GyB������8 ����:�=�g��;�J%��9����M�bc率�_�O���lx�S���\��Ռ���}Z�b���r��5l�p�m��-�Ky�&s?YASkS0�U�MB�,\nt�*&�O���v�%8B8�+�a%�z��(%4C�fVzHԃaM���"w*a���g�iΜ��Cp��ʊ��$�#�����2r�h)�}]�g~�(	kX�@��_#�h�x$�)J$c�ӎq�W���;�'��,�X~!�P�T�������.�d�>��N[�6`�L�x��b�?�tw�W�!n1���(�ȼc�E� v2ir�{[�1�VP�g���y�L���a�{��k��ݙ������f�F��3/�=T
o�L4��1$9z�B�*V&����J��aq�M���K#F��j3<�D��D���Ң3Vg�j�e>ݷ$W����"��]���X�
�c���UU�O��e���������+����d ��N�/a��
`�M�6a������v����K.�뮽֮�s�]v�e�,�au����N�F+����34��c�	�\g�2�D��>���E%8��Xs��H�R$�P&eT�(�0a��s���$�p�,GD��\qt{�F��9�_&xE������z��UV�+���<k��S8��)�h�:���x������I���%��C�׼˫��_�4i��o|�a�mo9���n���^4�Z%�$��<�(��[�ӄt�BeϞ�.���ݻϙ�/!kRO�:U
a۷�{�X�fB�` ���O9���|U�M�~b�;�,����/��?�	��������ۿ�P��:W�iE�'��_��{Ga~��`>��a������ $�:�7	#�@�0a�����C�����>�O�ap��R�F�t�O���b�/���/�������4_��<���Q~I��Z��f����svH/�ѐ)�e9~Q<�KГyE$�.?�����y�=L���h��הXfW�Dr�_�������q�f7XG&�`�1�xιK�`���,(	����D����dP<�a}��|��_����|��6[�2�ޫ���C/0�8�o��A>f_��W�G�jl�G�A���C~#���FA��sl���!H1b�zC��8B������26�xb`��Q���jܞw��]��1<��2V�[�B
8�>��b�b ��Xy����*��pe8%]��.�@(Z��Q!4�LrxYw���~���Z1�B<`�?��c��{��=z�MC@v�B��&��\	�,�'��y�΂z��q@��]��M��8v�8	��ɷ}��>7�a��a�7^tx`�Y� K�>�{����c,�'���W��N���$�	��JqOHR�s3��{�[��5{��������F�^@��З�2�H:����^~�y)Vۥ�dK�j֘��YO��͙s�}ꮻ���}��d�Ę�E�→
�����IfO�zx"8�����;�b��;r~���{P�{^�=`�{�P�OE!¨��p�������X��YU"�[h��^JN�o�rۄ�����(72.��%)h�6k�ꜩ3s慾/�k���3V�y^�8aq�F4@�BtN�]��J�QL�(]�s�Q���C6��0�1�ٻ� E|��y6�sƌ=J$u���hc��߁��T����U��5����Zd�����\GYf��9��g��{Bʁ�g�i���� �h����X'!��������+����/h�D��d�;k*a,,N���E|�c8��c��w_9P_	�j�є�����(P8B���y�ɑ�SV%�9*��������"�����F�W�q����
^��#���~���5��8$�[��M�u�]:��,���}T�����������������%;7�x����e�ƌt�N|�xV�\H�\g�g��1��a��4�8�p�;%�V,����0�i�UV��+؂�|��`qe��	���_{M�}u(5-�J�Z <������u`b|����7㇃�Q�\�0λ6�P��P}RRr���;��� �f���� )w�I``	ʕW\a�b hx(�/����Z��,1����2`0�u�E��m���`�"�D�,_x�E1�e:���F�,�����`�s�>gٹ�2�>n���iW���(^H����+Ì�2XzFp� (0L
�!T��T�#@i�C��e��C=�����[d�=%E�g2��`N��K���B0���lܸ�75s�+1�S��-!'�R�<������C�v%v��	�� ������o�����\��ͯ�^�w��]b�l����Ͱ��^e3d�q>�;h�>}�AY���3>1D1���a ^;b��h�'g�ƋA�/����C�Y�qǕ�e
���}�CPT���z��3킙�<,��j�]��V�^z�Ev=��	���_%H׸W��wP���P:\'/5�X�"�E�=x?~�j�G�O�܃��~�������w����y���]������:o�ys�
7:ɔ��O,�O�^%y<�MC�@�7��ЏF��iL�E���#��o~�[�BG��7l�qB)�X|��]���0`�q�{�Xu����؆�I��i�V7DP��B?���Dp�h�R�7Jˮ<�Yp6�qV"i�nͻ/�����a5�P�#sc%A��Z������?�A�d��n�y�U
(�+�RRI ���	�
�C�.�8]�b���&�5G� G���[�h}�Swه>�A͋��믵�g��J၄y�r�m�����ٴy�=����s�V+��������wER�4�U�P���̏l�'4wժn�����m6��̷WDC��AY>Rd�{�n�0��
+�8f�CZ�p�����MJm����ї�������6��+I-Ӂ���Q¡�����Þ,�}�))��Cz�{Gx�5����Z������]QC�|��e0��U�$$������Fo�x7�Ia1�i���9���haE�ߡ-� ^�Q�q�b^���v0xq-Y�ԏ��C_�!��>QY���v�()�y���J��8��}�� ��QI�=��Ș�c��^��̙D?���B)�UHB�w����-[}���k���v��#@�Ŀg�O^����q� m$�>ƾ���2'�J_�he��iq�o������o�)~��I�N��j�w�����go����BkA��D`�6'�v�r�ރ��� J�$.H�`��p��>� �G�����MvQd)+w���#H�����#�!1x�HW���Q��ٿ�%=!����q�z�-��8{H<���H�?���1�	oۿ/�ɣ�	�A��7V9_z�e_�d́��C�G,j����`�¡;q2�}�4μ�+VXUuȜ�J�����1�62�0<R���0��M����l�|�}Ùl��7�t�hI|Z<w�t�W^y��Ւ�/�3n�׾ֻ�Rz�Ӭ|��$aN��R�4��t��y'H秞~�$���
6�*+��j�3��p�uF�+��ǳE�� K�̼�ct]%s�:�4	��/�����7�~1NV'��](�;� �䀘l ��C0�V�;_��Kh�
��[N��֭[l���ؘ��"����������+)E�aNwe���/�	b����"�zԨ2;o���m�0KBw��@���H������j�����bv��0�:�l;[Fࢅ����ᒶ���KQ�핗^��>`cƍ���Lqoݾ×�i���F�9���S�7f
��H�" b�x	� =��'8{2d��Az߈�\0n޲��J	�eo,���M<ax�x�Sy�Ҋ
�l���zg��Y
1�o69-���>�X�4���G�H�G��H���:	�J �Y�67#8h$?��ƌ�}C�@	c�Ɣ)g���\���B��;�'ځFy}�7��I�,��O�����do��z�P&�aQ���VH�̆t<�3.8�rePSOҍ[n�ծ��*))2�r��1����^�]v��Q�b�~++�#ٰ~��pF
)99ѕ]o8���-{=����F	�iY�:{U�{�´E���ҁ� ]2�#4�	-Z��t��? S[��		tW&�F���*�a�"�g�\):�a��l�ୱ���SS��tT�`��=I t�D���^��i��̑�Z�w��=�Lo۱َ�Q�#͡@���熚`$u}߾���R�^z�u[��2p+��2Q���[<�
*�x�w����q��dY?�����*ai(>�Xo�A��J8�K����pj<I?|d�b~���)Fĺ�X1ee�~a��������k��|5�=p��⤢�57I)�8�%E�v��!�ӭ��#���t(����R_�6�/s�K��1��p��ŋ���gFQ\����4�81Xi��I��J+�s��PU(���Ϗ��/���x`�^� �}����קO��
c�#�<ao�~�BX}���k��]	e�IjH2��O��L(���س@�BV��/G��D>���b�-���L���^����P���.:�ϑ<ͷr���m���$�#dcm]��q�v�5�Hv�v'�0�8gΝ>�Wt/Z�wv��/�S
�p�d�Uj�dh�E�#����whޟ���VqQ�#��U)hY���S�!�%Q��}�{�}�w�w�I9��V;t��Uz�M�Y㖚��#*�%����x2���@�xv+��d�I��q�Qt����<حv�+�u�9�����Ի�.����ʸ��47y�n��\z��H����@qE��c�9*�����ز"L�:�,(��TY��j��v����1��~���r'#��9�L��@�����Dta����/`/�)sZ$AS��ڧ��n��z��b��o������vʔ��JwY��o|3R�[N��k �f�3���`)�s��(%o�ܹW����׎���b���V��,%�dL�r4n�x1�7�`R��Eb�Y.pXyB1���}�<�T1FV@�8��'e�/
̂8�d1S4J
���)IW�a\b"xa�$`��q��k��w�]��n��f1�<g�I(8��g|<�A�xȉ�G����E̚͵I	�[��q8f
�י6�O�e_%�b]__�{^�$`�0�w�vI�`8N?A̭���*���*�
N�l�fO͛�̓�1%��g뽬���L�x	���T�JB�G�3(݄����DJ2
3٥�=�hK�,�M��//+!$�$�M� � oOl4��R������<4*�����B�� �>�B	���x2��� <�SҼ��(D+EC(�֯m����&克�`A1b,)����9G#آ�mE��o_}1��ﳚ�4HoLX[[{��>�c�(�k6�3˖J��b�� ̜�k�H?��lG�,��E9cIq�*	
��w��1��2+3�ҥ��D�p�b,�J�"�w�}(�j�A��1g��{V2HC�
�r�d^CY�!`xg	��1�X��7�0�c�"�0�+Vp�Y���\8�%{�REd[�C�{��ZZ����C2L��_��p@��&�F�s�$���B�E>n�g����$��n�'��ǍJx��1���s��Eƭ�1cFy���l޼Ս�|�CV$��Q����
{�P���_��#VX]�6{�q�uH�`8�>Ɗ+4La�je�9���$���A�(��It��8p��������.��X�=�:@����B��G聄��#
5�ce����Yg����G��lT�?@/�O���A�R�<�&!�(�8.��T8�G�e3��s�vP
Y�$,��Ә`P�+�O`�)X��	ƓU7~c�G�>	nB���oVM�����y��ر\QW�\������b�I��$���/�akͭ��r��/N&�"�V�p ���Q�ه��#��;Vpdde�q�|d���9ٹ����M����.��8���n��f?3�W^����w� ���S�p���?N�4̻��	+�$R�h���K�&�2�����|�->�t�+�LR��H��_"����M�yY� �h"���#h���N�Nk�l�vq�`�
� .dI�x 4���d~� ��#��!�S��mgO9�#[�>�&k�1��)�dp�E�xM�����(f4%P�kK��x[�h�e���%��l���~0wY�bo)����:�+�K�%i��]f�<�ZgO2s��|��${�[2@pN��+�-��5��ǎ��[��v�{�i_z�Ӭ�}���=z��Z_AB)�lΥ�a�l��y�YH��@��`��Q���U�4+N�_�yO�6�cz�j pa@�:�X�h���aE����=;��Jx!�ך��`�ѡ��d�P��Ha�0.�q/�H����r���%��=�y�tcc�kڴs�a<HQB�0�=�C��TX�}�=a#GW��l�62���6LI����:"
���ECN�4^��g�0�R��]�"0P,�� �ҷ��F٠�C��b���EБ)
�
�$��U-�+�:E+M=�|�����Y�i��D��q��o�`5c֬���E�� ��o/�p���p���| B�VD��v�I�N���<�/��սD%'�� ��Lwo_qq���B�r����ـ�2�y-����_�Ņ�9���F��j[%%e��Q6|�p���kw�|��;>�(=Qi��#�N�'�X��|����,\�����^D�=�`@� }��q>|��B��c��E��:��a�Q�N��U�6\�l9L��[2�XI�p%�zb���t��[�a�Ђ��.V����7O,<㊢��V�� C�4�R_�E٫�8�>�!��	��8v��:���Y}`�U��G�=\��v��1��~�1J	xe��1�`à#L�@h��HS^�s�s��j5��5o�qxHJ7�� ��t/�{�!"v��ϱ�1��/��*#�{M�w$��������
b1���?F?�j0�؛oa��駞��S��`��;\q�jƆ9�kH(�=$))���j���T���b���%t���l��R�C�+NM��N�N#xf��0+�d�|��ٗ�&�a��;w����ӳ�	&�N�<�������`�0�ǒB���ݻ�����?� ��G0����E�<o��}�|����,ɝ4��� �l�AH.������wPj1�����^X�Ei�i��k�z�Pc�Y`^0���ܳj�aD��ŲR�j	N#JB!�g�@���-a��i�@���'ΪB����@�D���W�ɚU�l��;�B���,���n`��������?l�� U����cL�c�c���yl�K�nIQpz��+v��@�ц��wCn�9@��K/���>Ϟ���Wi��\�󅬜���F���bq�9��(��'��K	�'lʛ{�\��9F��#����HT�	�UI��` #˖/_髣Dhp���	�#�*�V,������8���Ra��%ʠ�

rŗq���[>��h,�[d'�1Y��+c��@?Y�f�'�y�ŗ4W���$�� X�;�����vɬ*O�t͵s5V9��t�+���::Z*$��Q���_��b�N)��iV�듃�,].�t ��L�+.�����K�'��g�ּi%}�%�ɞ�!`����'SJ?JuUM��O/]�CX���
�I��#e������XeH����I�>k���(��#	Ɓ�B)��Á1Do��L%W��+L~�a�(6���]�Ї>�����]oC�qfL;pab�anx�	'z��'l��v��J����Eˌ����,5��` !t��%)�Z�{jI��t�M��P���, �-fØ���9%��0+��y��j7x0�p�������n ���R	���#U�����@��0�a������o���ᖛoq��`��[|��9R��%H�� 3^�eHA�[+���!�qB)""1�
B�x"�ߩ
0�����tO$]:�X�����yR��P��ز����1��<-��d�"�N�z�o�f�{�0�Z(���K�٦M�]Qypz�,(�:q�6��~ȨW]Y/Z��u��2���{0dp"��=X�Ξ}���5~�x;&c�M������\��BG����4�2>X!LF�HibuO5tF8
�IwMm��B_���e�`��O�l�27`?��Ox��9��6LF
a^�#���J^�@���7��Ns2�gė>�2�]���lijp�(�i1�zE�?�y��G}� g��{V�>�я����b�!���,_R�QQ����#h��Ǭ�t�X"�F��ƞ=#�D/�=ι!�Ŗm��3�+��� ��	�a�b�18`�y��4�?����o}�Wzƍ� ��,�'�(��G,a�-��$��`k�P���OV�*�˥X�Ә�����Lg�j�ax�-0%-ɕu{Mop�܃ga��nQpq*�V�}U\�� z?s�9���¸�ڍT�ȨTz�9)�!�CV��Ӵ��&�}e$����������#q���9P���!�$�PO*I~O�xECc���Ck�OV�(�8|��xBY�݌c�NW�u��@���|!��MH"�[�#X�fHY��i�F�1��LKO��v�K8����FUaq���q'4��}�7�p�U��̸��?,I��9����������c��$=�y�3T_處����Z���8A�-V~��W��	�ʳ�WW�%���xRpN>���f�&��R{��D5z�pkV���	�%���c�7A�s)Dk${Ҍsϝ!k��RV�1B�c�J%��PLx��87eÉ��c���=<zc�I�0���]~c��7���|�7��|�Ig���<�AUu��70�|!҂���x�H����1�@�,,�Σ�>f����m���^�z�<K�,7�����2���+|�=99C�"�V�\�yhG.�p�㥥7��_��Ho9�K��t�)����/��(����z���^#<�'�=�����,�Wj�Y-ARUu��Z4�a��BY�$�Cb:����XQ�P^=�KZ~ƌ��[��9oƹ�IG�b/����@�"l`a%�?)\�`liI�T���k�9�%�L���dg���n���lD���S �P��I�Ώ}XW[�����9�����`@��W�z�+�b�20��Cƪ+������٢���+ʁ�d!"�V�`=�����|�ŗH�ɔ2ر�� ƫt��1F�w�S���o�A��c�+��=����G��b�j
��(�xk�͟��+x���/���G��N�Fa���]{gP�1��3������.�h��w"��Da�'�YSS�6[]C����;�D�2Џ��V���բ1cF�p)cW]=�ƌ�J��:��6K�L�q�g}�ÁR�F�E����Ç����w�!0\���` �GX#c���E�T�=Y�Ҭ���q�+]ڂ����E����b/��%89�<�=g���������l�rw@���G��4{�/B����R;d@HP��_�\�y¦�T���al�e���}
<I�yR"��9����>�<���M�2��]k�0Y�����81���w�����gkK��L}���aC\�"�9�?�:�#
�Ηb�7��;��Ǝsb��"��\gL��ᾛ6�4w�4a���o��p���K�\�G?��Ą���d��Kr����8o��U
_�Ӣ��0�J8#pJ��t��`/��+�ۗ��eWb��7]|n��a�(`q%$�;�W�_w	<���1�ۭ� '���:[��x����QP�<�>��ǍgŅ���m%�=n΍i�o��RؠSR�C�|gU'������2(O�"�X�g��G?z��԰�	g ����-֘q���3��J�����A{\��٣����� s��@�{A�vȼ�#��g�+��6�5�j뤄�Qs��8W��0���U���Ɨ=�j�WpN�
V��}��@ '����س	g8���q�Gh�S˧�fh�d%���
�%E����p)#�d��i�5g���H�rF�@����� Y���a��n8p(ifF�Xb�^{�*�����_����83�Hp��4���q&8��P�FqL���M�4�N}!����z����ƙ���t�R�O�2��#����]�p�mܰMrx���?a���#��%Kް��*�DΉq<�xBm|S�ˇI�X�Vs�ʝQw��"Y����*�v�'b�YNX'�*1�ެ�c�0ő��y�@2?�)�3���s��dN���+."�E��_+�D�Ɛ���,'�(!/�{�\��Q&�N��{����!���y�Ә��QȚ�@_O�_r9I:I;�����|Ds��~�l��׿����ӿ�H�Y���>Wz�������3�M��Lb����$A<o�S�v�)x%�uGIiok�c���ns�YR��H��.�J�5�GK����}֙vδ��Ӥq(��P2{�2�����c�OJG�34)��#��X`�0�����QE��geU�+>cƖ�i����t	�fk�o���&k���/��]m�RĆG� `z���Ce��eRЏHP_�iz��lϞ���[J>o�v�@YupPx�S��8DQ�+x�Q�<�,;j�ޝ$�$x��!�V��5��%g��0%L�/ួ{=��G�7mv/���\a��zPj���|�Q��M���w�O��`�)Ϭ����
��Q�ƴu�6�Cp��#)��V�@�b|Tj싊,=3M��r[�t�p�O�"�>��ގxY�.m�>	n�B���`������ܾ�7iO?g�M�0N�+Y�*5F2Dj܃�#,]�c��ム~A+��Ч}{wI q">���{�u�%�e��DA�s����%A���7V��+�l��2U6���������?������׸�5'�r�F�=�7۾����$$c g�Q�S z׋��q��\�H������j7�&O�dC4��4��j�e��@*)R�3]8_#EO��9�p�}��~�i�j����R"���RH�bzz��7�V��QW	�	gCNRd0��6y��cg+,�s����A�7;�2�x�g�8��F�P�i�Q� Rs!-=��'�m�xI��u���%M
�K��l�������F�q+�2�8����:~��`pX*��}u����C���IgH�!;f�{�	��0�;g�`Ȯ�$>'BQ/��RM�[��u_�� ��_(�'+�a<����/88�����!�J�4�B-x��7<�ٖ���jA�M��s"췃��[<�[�����IY-(�u����5Q�O�3���|��;��d�i ���bC��r/-�yQ�Qx��^�_����ij)��W*´7�c�|AY}� )@ֿ�ܰDq��)��E�S�	�
�|N
V�"Bo��z���OI��a����Q����t�@Q�ޮ���q�W�7X<�}mG��1������b0�X�d��F|;�Wr)���2�<��,~���Q��բ9@TA�d��6�⋥<��a�����R�ۑ#ˬ����B���J]��g	N� U�$�f��+ˬ���翰�[I�/���C$��3���j!��9��s�M󰣽ō�jA-M��lߞ�v��B��K�u�E�J�������5b��¹��e�#�=��W^��
8����k#�����&!��2�Cs�pڑ#�Y���O[et��;e�Jf�+@!M#�=&9I8p��{�>25��|���=��S�WX���X�+D>�N�����Z���"�WP\�_d���&�ƛ$w:}c�s��+��Ƕ�k�����dPU	g��+��>3�'�@��Y�}�=H}��D7��ii�&�=��㒵�Ǐ~��t�֯��]�-�u��r{�iQ>������t�����c�i�99�g�ޞ{�|32^R�#����-rO5B�}+C���'H��Vcg�9٦M;W
�()��c�'�}>.^�?<a�vn������G.@�qF��r�w��ChcQ#c��(s	�(B�bVb�G:\J�٨Q#\�hM��	$Eزy��s��P�+i(l(&5��d�By���
������;v�p����:tF�E�A��J�+���N���C�x�s�n��W��;�����+����z(�w��P�(�����H�����a�A}����?�T�k%�
+N�W����h��D+�r=f�X�Bb�o���׋�x��+��2V|b�nٺI4�g�b�J*+ba����0(������%n]�#!ah�w��ӥ���>��t<������X�;�2��z�T4)U2��l��#I.�,Y��i�$CϹӑ������h���^W���1��I ��g����?���m�~��:��}�n�l��-�r�"	�r��-���^}�5�:F���0���l�����(�\c���zD�l�|�{		���>� &G?�y��n̨��h�rP���k/�v	u,���V�b���YY�I�3�](|�,m�9�QR�ՏcRXH�2a�8��O�F�xC��!?������%���m�=>7���K���
��]:,���O/�B�p��/�g��Y�3���ǟ�a��@�����Q�"_�XtW ^U E4�{�������wF���n��3ha@�{�)[�v���|�C
��+��_�����gHR$Im_-4�xn���ں
��$�Q�JzKS8���k��bT��1`�c�*����l�햓�����uG�7`����u�s �8 0PJ�;��h��>�K��|�]w�վ�>i�I�C�YA&L�UMλ������|�5� �s�q�4Y�֣`u�B�L�V)���������~��{-'+����� E9;�U�_	��`H�b���w�`�Lf��5�<ÜH ���l�
��A�;�
�&��O�G�����f? Reu�xhXyb���2�F:�@�����QP��S�Sa\	Y+-�+%_�����q��%]F��Z��o7���N���O��q�M��J�7�`d� ���178̜����K=L��p��X/����+�M���?��x��t�j�3�M��T���?"��Z=�[��/-��ڈ��6a�D���>n�X�#���Ycw'�$��ē/�}�}��{~�gpd����]#��L���'(�h�.WTg��d��� �B�;~�!�9�7����$쭣bG&[�0ܩ��ֽ;��UU��8	<�Et��V%}��.��B��τt;,��G� |4֜y�EC�����+,��Ӿ�H�Y�瞻�VTT\|�رax��P�Ŏ0f>^$�*�툰�FV�&{f�� q.� C�����L�|�8P�m��)I�v#��'{�]�j�J�F����ҿ��i6���ҳ*C0.>��Xt�}��p 7)÷o�ឪ!��ٹ2��^u��Oe߁}����٠CC���BxY���J?����72(�T{��pR�>)���0e��p�5�Y��f� �S�	!�'\`��/dS*<@;S�H����lFV/1���i�g��>2��_Z��QE���)���(ĝsH/T�`
�hBP �j"8Qv�ۢŋ�W����� ahDACu�Vc����[�k'H�p�*ly�mfJp��;�C;�<�_=�����gK�
����FC�=��cFF�M~��B�UB������%��?�O����b�wJ �ۻS�N��	ƺ�6�l�{v'Ng�F�C
�ue�Ūk���E��C��W	����{���=��4�� A��� z�o���O.8�1��n�n��� ��X/!c!�g��Faq��\&��I�^���f[����s��y�o
�Ţg��L�"ʎ�N���Khc����!(
(𬄲i����aU�T�b��	�8�9g�3}�Ka>Q�����JbVk��G���$��n�;~����7���O���N}dXr��h�(���C��Hiy�8od��u�m�f{�g��{j��+���p�g��*�E��;�_�`$ A'L��R�� oX��c�k�#��h��|H���B8Z��	�'~��烱�Exan�#��7�a������_{��c#��)�{�[ga<��8?��ٓ»�[�3����>��{|3�#��As���G�#��ʬ��<��>�;)+ҼZ�:�i�9�J	��歌����5s�]v�e�`�|{��gD�͂�Fs'Q�DX!��ÊY��N�\�?(�5���F��I�x�	_�`ԝ;w3�<܉q����A_S��i^_$D��S�ż���q�r�\���Ϟ��.�o��7��0���U�h�����X5c�p�	~ �A�����S"yN���^:�R�0n��ڴ)gYAa��!�GC�m�Mv\��*��|Æ��ʫ�x�1�f�#�َ���D���g\��Td4d��e�w|�3��^f�G�����@R��.+�60Tt�q�R&�n߱Ӿ��/ٯ����2Ńu�1���`������'$U㌣���ғm&�ҨQaU�� @������[ 2}���p�˞{�E[�x�;���-Ex��*��l�lJK���t��~�>4�O�~��#Ƭ��׾ٛ��Rz�Ӭ�u�'�J0��$&���D%�.?�H�E��g���VB*KBv��DYf�*ٜ/Y�i!ܶu�{�P"X�߱}��ڹ�/Zh�������}��W��P,XRB�M�<���T�N`N�)ug�|�Y𾤎��a�W2��ɖ�e�V�

J�~�)ǘB1�8a�z՚u��C!���ْ%K�1��8.���S����y!b�@�K'Ư�2���u�p9�3�w��}���9h��Ͷk�.{s՛��˯8l���r�B�A���z/���_)<���^x?w����+#���
%t	#g���M9bK�-�����>��wl�pE��B�@@�_��7A�G�Z�M"���,�&���()��-Y�4��S�a�+���}��R�y�&[��[-�r޼yv�}�������������XzH���� e�B������R�jl	Ôbտ�8���%`9|�����^�R
ܓ��el٬��S��cSN�'�/2Q��j��.�3�(8�_2�PzI�\.���%�k T��x�Av����R����J�����/�h�-�}8k׮�yZPX�khjt�wA;�P��ɻ���i�p��,��Y+�=������Y���,�5�~�d)c�1���d�R�����ɢ���,�y_5+cWBG��^Y_%�7��e�$+]�4�xb����j�{�{��$[�ѳ�=�F�+R����ч��;1��ο�A@�;�]�r׮���gAߒ~�+�5?g_|�`h#G�8WȨ�*\�%s���h\q����_VWp��u�0N>l�� 3b��g?��"M�(����6hN�pco=���_�����ϰ3&���{Vŉb`���0�����h(�
� ̎G�H Ysc��)����~�8o�LI(����9RD'N��g�<�@fY3|/� P-�7�^�?�0�Pg�dV�5:�_� ��%≰���8��%��Vtf$�	XYY�"=�۷H<:��������'���͝ns�?��"O��xF��HS�aN�K�x�:�(���v(�ƃ�&�1�j*+d��[J��OJ�"0�~�[��\��V�]m�/�o�=��m�8���J|����/al~�#T1ǥ�4�՜e����TTT�A;v�x(�g���o�n�F�'r��]W����Iz���-W�6�xk����O>���+�A�l7��R~���f�a$��ʫ쬳��!d��n����	�c<��C��_�V%�K�:|�����$�̸W]}�w))2��������X;{�E�_{��YV��w����g����������|��DK��Р��?4�Q+�Q+"���*�G�T)Z��-ZT�CT�d��Lϣg���}���g����MԔ�T~���s~����k���Zk��������׿��BS��I����{^���鮻�������K�w�����o~A=�F��������=���/����W4���,
`~��H"^�ݝj��;*��;[�����,��f=tm�����e�hc\lfp��Dp�@m�����T\����ٳq��o��zhh/���ԩ�k�b)�I4���/�[/�����㟬��٦�������y��UJsh���h��i�G�o[V�X��}^�Gj����͔؅̒t)wva�"L"���{	�c����#6�iuǋ*?�� m���@:��I���Qbi%�p\}5GqXΉ�Қ-:���cxy� -�n<��9%����3�XbW�Ƥ�]��2��b�2ew�3`ے!�e��9��ό���qu���ȵ�Z��@m�zXβ����ֆ�_���!��%o����m�����#;��|��=���w`,_��%�����rʼ�q�♚1�l�{�Q�>������n�M�.Ýp"$6�gf<+�tk+t�=����EЭ����Ͽep��[���>䫷���?�v��]�`��1��k�����Vږ�_����� =m
mW�01�.���pd�����X��� 3R"������y�[.s�P�E�.Z}Ѭ=�Q�m�b�G����}<K�MbXtVx���E/��kw�ѝ����e/��e_�ڨ�N���Z�g���~���6θ��in7��tMd��#$��&��\�#�����i\Hz�$k��j���"�Ͽ�c/Nޅ��8M���rL���A�o����x��`ck��5f��#e�c�{�
��IޡEТߘ����_ҨGs��{I�����n�5<{qtš��/����e_lڪ����؏��f?�#fȣ<�Ufoc}��
�"M�n��(	"R|l�n����j��B��A��}�DG�����y���/}i�hK5�(�S?�S�����5�K����M����h���}��ކ]�zZ�Ƚ��$���R3ާ�YK��(��E�Ɓ�?�:����>b�#�K�����R2��v�Ccцg���&��^���R���/g�gΩ��yK��[/�a�������.�D���#�����|��6�/zo��z�N�-Y^Fw�ej����x�����Qґ��G?-/V0�^��?*�9��S��5�X���wٚ3ߟ�X�˿�˃�|�{j<���6e��e$:��}�m�Q�K��K��<�}>}tc0�o8��g���e_���s9�������ߨ���6Kj<�o�7�/�0c���=x�+�r�?���7F����<��o���Ł����������W����S=�)\��K��N���?/�G�?��~�g~f�A��~�gj�� ����������wn�����g?��QBQ&�))J�ڷ�ˋ+�Lh�I#��\��1��G�X�Y�|>�)��O�!*]ɡ(*�r)	
M�f�<s?�F:��p����"�X�(�^H��e�r�(���?rM�ȩ1� j�|�q��@]��r]��p�� ��d3^[�.��/z��!���~��Z��=:��97d�i̍�����'>Y������ވ1>���;-hP�{������v���pY�A�S�j��=àHi��r��&��\�K[ji��o^0�-��1���l���ld���+�׆m�7'��ד�Y6TQ�ی�Jn��!����f9��P ��ŚB��=��$t^jK��l!K��5:����y!r��=$7x&��N��ᫎV�m�?z�H���Qn����{L}Ý��̀���%/�p:ڀY���o��5���d|10��W�bee����\��g@�����g���"��3
.��ڊ�Y��2v����
/S7���f�ʸ�o�ٍ��i�_��Ơ�|�Z�3gAS�y���ؖ֜mzC;�K�Rm�����&���c���E�o�Ѯ���Y�)���� ��p�δ�HK���n�PrLl�������'��<b����o���R��M���[���{~�|���R�j��-�.�w{���s)�bOA��/��7��v��NC��d�q�q��c�@��C3X�%�q�w�&y��z�u/�ې�Nz�������i�ӑ��ڰ�7���c����r.���L��>�'�����`�����ޖ��C7^]�?����3��>a �_���h����	.p�}�w���]�E�y�n'��즥��q�ɪm����n��v�m:�v�@��碑��B�����̾�":bR}����vb���_��5�F�9S��A��>P%��5���f�j������_іkx�	J�B{��5iq~o�C����C66J��];�
B����O�7�W��ɇ?:8}�t��R��q��"VLp(ZЧ�P��-	v�W�Ky�q&����{7Q������囆/z��Ֆ�*<C��|���[��[���,�_uU���+���$o8o��9�Ԯ��>VI�Yr�~i��t��;�W��[����љ�n��`�`�Ȯzx�_��-��_��ng�㠋<~����U�_x������������۾��=z��[�������U�:H���M�J�O}������}�G��mo{�5��O��G�{,���^��?:��_���i����i5#C�)~���� `�{����u�Rx9,c�{�(�A��S��a�+�%"�ڠ�����F�o�(��d�(Ϡw 
�)\�z��u����3��N�vK���L�톗���]h[�*K��2��l6Zi��ѓ(Z)|߮X^�;���{J�y�� mC������g��2+֖�1^���e���l�&墥�G:M�Qi��|���tρ\����f@4�8#A;����fD���`Ԗ�̭6sy��1
o<�dĈ��VV |��I��V`�ᔴ�Y���%"�������qX�f�p���h� Փ'_:��9d��ycSM[RK��l��e
}dk;�.�@�{�;�'�k�]��/�ۮ�V�ޕ���0\�摧�t�v���۶���jC�#M$��O�� Z�wXe�Q��⵶�Д�3����Ň��~M�÷�1�������Q�����K已�a34l��C�s�4�x���<5C�odm��QwNt[�exeW�!?>6^����%�9�F�-|��&s��3ˍq~��=���uM��\�G��m��=-��rm	S�'2��X�]�S�E�'`���]�4oO�̘5{`g�z�#���,��I��^����؇�h����v��qP��9���BC�5���Nh��@��!.P��_];_<��8��۶����<��Pe|k':��1 A��O3f������-�ɞ��m�iz��0�̶~b��ͪ���GpM�9�O3�� }wm�G��Us��l����.�t��Z�4Y�fi.uʽ
@Dj�΋���B�)��9z��@��s�	y3�����=|����Ap�}��[�� -��4+��ÙȬe��x�	�䏄
շ�B���J�������Sp�z}��fT�3�nk���`-��ګ;�p��*X�S��fm�����Ƒ��}��?�E�~�$�q��m�ku��xp��ɺ/�U���xS�7E^j� ��{Mg�K$���WBv�̷��m���y'8�y6�C^V���V��E����MNjk�N:z_����w��_��_|�φ77'����~�7���jp��#��g�?�����4�Mኇ�a�p��C}��Ǐ�����ַ��������7�K��O���yv��w������������uޱ�k�r�J�+��t���68�E�E��+��z�E�$7�y��E0)����
�����˨D�����h଍R6%�`4�A��u/��6����	>� ��8��G�>P��r�|���)�f��M=;��NDv�:�D3
��p�������c �-���;��Mz��bZ�h���oD����z~\^���Ð��`(��׍�nL*_�:�=��h�����-��?ڡ��5r��O��A��(��$��Rꇝ�T�c��(�gQ<+��a��+e�1�Z z��{^�-��IF�?x�q���x%��4U�'����ȩ�L	:۸ӌ0�۠]�߸�w���$�3v�[_��F�O�~q)�F.RCR&z������-���8�d</��^��<�-��:����(�"��h�}KB���x��]_(���Q{`(Y�=�V3�`��Q88�嫶eIfg[����K�9O�1���vjF�
�c��Q����Ж%7�+)J��]�$Iy�l|�>�O=b�/x�t�?P�g[��N���sX<�Q�Y���ǎ^�+y5�l�';k�6SS�W�)�<�!r�}��h�N<�%��/�_���66��e6'S���3=�rf�'�����Ϟ��;yh�N�4���'>{7H�q�� t�ۭ�^0�z����F/��A��<�b�t�z��1m���>�r�~A�:��G��M���j�����?��T2��f/�������*��[��ڎ�cV����vY�Vx��0�`������lIWK�f#�8�S�kyz]�-�p��Ȉ28:�p��G�r�'gi�fՓ�--�*ۧ+|�)IJ/��fm++Z�M]��N��J<�i���M�j)p�&ޢ�n��~����^�<~���jh�	�ێ��/#'m�mε��	_\��tB���JN��j���?:�گ������΁��׽����;�[KN��O?��bd}Lzc{�d�&	���oڌ"%���Nm��x��Y�ш�����#�=�e0T_�?�K�
�%�ک��`���E�9=�'zo��`�?��>p�>~�]�W|ٗ��?=���S����˯��^'l������+_������9�+��3�+N�xp�ɓ'����������-/�"Z��xSE�y���'�����~�j+XJ\Ǿ�Bv:����d��"��(�(��(	J�`川Τ�Jet52��+����Ep���� ��y�.UJ��_�.�4�ƒʪd��:�h�å��ͫ4��J�C{��,m)��Q��(�(G��K��ً�y�=�@1�� 6W�,;q�=s.��%�{6K�+�M���hp���1`ڌ�¢6`P�FيfS��n1�C+灓�K)j�u��a���[/6�x�0J�=o���R���%��;'�ޣ�-���˓�Kz�yy�p�C���q~�� 0�p��P�ީJ��:31��yQ��1@˘H��e�ڍ�����(�@,=Zi%��� A]8�]��ﴫ�~��I���}E3�=�c��x��}�8��E�����b`�X�ٖ��	J�Q2z�o�i_�(�����?��{N��p�\��3�Y��)�E���'ksI���/�3��:�?�}��;Z���G�q���or��͸�9i?�ȑ�e]5����%��h�~���/mɇ.4��2�mdD�A��Ҡ�9���xӌ�f(�ڜ�`$Y�葹���vt�E�l�uX��t�Ѩ6MnZ �,Ԭ�H���4yv-�.�^���5�����_:#���^U'(|��7��w��)�T��Iޒ��!<�M�������_���a����=�;?x�`��5�m��㏷���T�t�g����ѓC�ge�ŹM�ҽ�<u��-M��tB��B��Գ9jq��ԁ��n�6� ��YI��<� ��3:��	Α�)m�v7��f���Z����qɶ���񔁿�ï��F���G���ٸ,g��.^������{���wms�p�g�/RG|����-�ܜ�¥�/	4�hR��?2c7J���Yst/GN/�oc�6��U4�x�ءh}�*����^��̆X)��=�������U�)�/ڱ�85�$m�Ggo�r�V+qNl&�=�B@S�����K6Svm�9%�vƽp��K����[c�w~����苾x��w���Y�>R�J~����ښ����K�/����-���-����bz�lb�:��p��y��598H5�������9��weA�������	{��9Y]v�ݣV�Oz�=Ws�,���}t��_���{���s�A2;�������7�	�p�?�����kߕ:5������0��'?q��?����7��G�=�7��>���/E��}�<����wl��%XJ�#����1������Z4���T�]�[E��x�d)��$E1��z��x9�׌4�P��K�M��֠n���q (!�gd/�� �>&ECSD/�R�f���=
ϼ�`�;��0�ш�Rh����S7��G;���� ��A���}��T���o�Dhf0�j�R����88}���~��=��C�%��ے�e�p����84����i�%��Eی3lm�c�2�'0jj�W� T�z�Bч�v����\I�r���A͵�bf+�cp�����3�+��Z~�-�>(y.tVd���|�6��X�d���vVjF/�R��n�9�2� ���1
���x�{F�z�)�s��qt�pHן���4����3�좣�!������w��!0�c��v��n�F��qn�c�5��z��Ez}7���ad0L�����}x��PF�xi���Ԭc`L���A]��b$�Ϡ���U�rx�\r��͘#7��KA� �������Z�y�'>i�񓢝3U�5d*}~�oU�-W�#���Y��w�w+��iF��7�V=��Pn2�[+����#ry��/y>Ih���Su˳r��������M�ԝ1�y@hE��nmٌ��^����`�w�"��[@~}^9�9���ImV���xGm+L^��o�?�շ�����o�]�|��SǏ'}듍��Rk��~�Q}�U�VK��cQ��%�׌�B&g�5�Q~�x��Q��t�^<{���d�����'!%W��Vh���tu��Zf���lmV�Ⴛթ�$�o&�|�gE�|)W:�ʥ~P�ji��Μ=��e}\���ܴ�|mV\3�P����~j��W˯�v9�k�B�ߘX�S���S��.~�g���rL��"O�,��t�s�Ș�ʂ���#�.�u9s����unN��Q��A2J�����G�;�H�?�?:Xc��~��[n���������O֒}��C9e*�>}����X�Q��kߟ�c	G�R��8��D:�Z�Um$���*h�����.�KzV�`sx����
��Z4��fwӦލ������p��3�p��-M?�-����_�������S��?��[~�ʠ���{������}gڬ��p gS����GN\}�]w���nz�O��������:�mn)9��(2��|��I�h?��l�VX&#���H�A�)�&FY�1����RQej��`E�Xnҗ���o 6������+6�(J��Dꪎ�<�T��s68)K9ͨm�(%�fq���'=ZY��ԕbl/��� �LE}�Ț��Uy.����c>��[y� ��}�2�����,|GGSyK�@_�H9l�~���rLmN!:ˀ�{��3jl�k�#�;�J#�/p��miG���/g�����*�.NM��2��{/f9HՆ��V;�":�}��?j1C�ݬ��=g���Dm�{�����ㄊ��À��6�qL���	���zs<�#�ڵ9v�k�^=������G���S��H�E�ɛ���C�L�/��%oiC��=�!��2��x���N�߾��xR<�O^��t���1Nfh�41��~��%�䶷m3��������V��?�U~7"0���|9�sg�V5h2䐯�����<�[���͸���O�Z��ӧ�u�>�m��f4rZ����i�?^������q�^.�������+����:�а�eØ�3�f���2.����R������{�RW�G>��mO;��۬ʎNV���%Kms�U"}��k��m,�|W���]_0���To�)���  S�P3t�z��h�k�Ǥ�i���w��/c+3�����9wY�mf���WՌ�t��S�0�^��8�t
�A�z��.�����{��F�2��m2��?���&vf{�/��G�x�'Ν��3&t�ծ�q��гځ���|�O���d�)d]�w�
��Ֆ���}6�4�U��G����\c�`� ���I_(G���On�X�O��:xh����Re��Z`t#e�=���2G[e���_})�vr6��,�/�����K}�V��և�ԩlr�aj~H�P���q�c_>	�\��WNRs�{�����#�ǹZ���-rUcP����.��Riur\r �bxm��M�<��Wmt�������|�w'g�����ʯy���ymDNኇ&�S���̙S�w�}��~,�wϞۿ�~�l�m����R��a�cfXll�����'
a!��Xc<|fq�(��8P�(
�\rQt.)�� ��(���ua;x8r�O=:fӁIP9&����O��XgK1��@Ӷ5QG��I�D��s�����(�I�4�p�xTK+£�-���ٵ�Sa}kwp*���g�7�x���Ϻ�)���7E��b-���Ȁ�w��u�����	���
<M�b��{y
�9y�oF��.��]�C����r�����oO��A����a>�����ԕ���c�N?Tb{����U�\�c�u7����;�C�-��'��'�����y��э[ϛ�����ǅ�=p����@���/�8!!��}eד���C��2"?#ƪ�ޓ<��ɺg�V9�zY?��IYΎ��˽^F�E�--�w�Գ��3A�1�^9e��|�'骍#�ڋ�_�J��.�`\��+�N^�����������n {��ަ��錯x�����mva�e5��@�}A���j�܆58u�'S�V/t[������3 �C��̱�A$r�����;ups�l �{�P7�2����=��D0O<3+���R�9e�r�s�wbwg�S�mv��ׄg�qt��W����~8�}'���6���s$�z�Im�)���L<�6BT�ԫ�g}�{.Nqi�z�]���s�Җ@���r�ա�\�
P�U)�@�/|���J?7�v�س��{�{�����g?�C?��/}���߸=�g�{��4���>r�;�����׼��/z����DltNQC
��AE!��跥��Ωc�G��t�"�;T����['�y��o�f�W��(���
��5�+z�ճ\+���96�j�:1sπ�� �e����Ζ����Ν�Ș(c��ʑ��Sj���S*m΢���:�fX�18�����C'��Oz��<��<����fW��_�p�
t������.ZD��mi��l�x���3S����i�m�H%^ Q����K�yM�Z/l�?�Rf�/�{d�_YR�ٳZG�%5��0�r��&y��L�k�1>z[9�%�v��yҟ;��m�}@.\���߽iշ��4tp����pO�d�=g�J7�t<���z���i{��s��ԑ�ڸ�5H[>v�`��d4.r��9�����Wݨ�:��
��e�oZ���>/ۧ�ʐ�O�.��+M�&�6���Ó����&� �Z ��6}��u��˪�D}?�G��>M7��6�S�I��@�2j'�蜧��g-oޮ%�f4�* ��9B������q�T�IύkO!%���`~��=	��V�<}�9��\�>s٪�06��q���ڌ��7�'>'�:+�y�L���#�\��<��e���y�+j���I�_��߮��~[�l�n6�l��w~�ǩwc����W��n��%(SxF����)\!p���Gϟ?�����/�Q��(����D!H�\��K���h�(��M�;�p�t�2�s�CS씌A�oʀ����9��_�q�o�(L�)8�Uㄹ��Z)[dN�?e�cw�����(�a���x��Fɣ۽�����S�n����sE基�r��z�#���%�L�mG��={v�=w��Ѱae1�h{k.��Bh�iJ�9h���=��?^&����=��N��t�Ms�]w�Qv���s�);|]��ͭ��;�y�S;O<��ΡC�����R��:��p��,e�x��Zx���<gO꾨�>���� >w��z����7��sG�:�?pp��C�v����M�x<LY��	Wf�F�kF���8_��2ʽ����s���~1�O������͍͙(���lvggs�������x��a�,�9���g����;ڙ�����g�b�[mv6e�嘍!1�0��gq���0����Q���f��md ��z�=22��i �#iFi�!�!�q�cge����v�M=�r̦>�9d��<��)=d��g^�!���9t��j,ys?Ť k#����%g��k˯�Cp�̹��E˘�qT�I#%Oj���Y?�-j	<�&��.c���'v<0��[_X}o;(G]�q�{�<��i%��`L���8p���OD�s�����;mw)o?����>f�����v<��^V/��S<������Ɛ�'��s[������ O/or���ˡ:m@rWx�w��G����g��R� ��OB�w)ݸn�^g�0������`��%�ߵ� F =�evd��#ܖ���r���~����e���C��G�8z>ti��4�]���Ug��@�s9���|�t�f�y�Mε�/4q����Y4�lL����Ӄo��+���S�~�$�o�u����&O��_?Y'���9)��~ϟ��������k�sƕZ����:���{��#��;C�����5��~k��t@>��N�����+�R߉�L��s����]W|fS�QOG��P��|u=��܅���3C�k�F.��MAJK�=x$�%p�ă�����}��ߋ�/y����N��'N�
��������ۗ�}8�������B�1{u��n�Ѹ�"Q`)FV��Ll���p{k1Ja3�(��]J��Z�e�ڞI'�s2�����I��<�H�3f�vn��/�wV81����j�]e���ɿ�k���VG踘�r��y'�9M43����0�	��1����̃Iʸ>��wBjeG2��,#y.ǁ�2�%�(�.U�߲���#*Z��S�,&�E�	[4�����n���\�n�h]ɠt(����WF��ʞ��������в/�bl̇��1�1�Ng`xlqiq)�o�q(�9��k1x����h�l|��Q�qPv��6�+!��x���A���ٔ�a���%:�]��p�f��b{�lFHR��Jpͅ�3��Pͽ�{oP'+e{{g8�3�37;��pf~g8\FIx�>;7��n��G˩˾�'_��Ӿ�[f�,/��Z^ܳy��1y��,����~�sf�z+���j꿚�f���B5�?���u;�vҺT�8�3�%.���ʙK�����U�j��F�=ɷ�4�I�$Q�@Jf/�l���N(�r�z
��w�'�쒫�3s����K)b&��d�M駣�Ͱ_�r̆wC��c�.����0|]��|;�����WG��s�� �C��F��Vh)�\28���)����׃c7χ������Q����KT���&�i����g9<t�F3'x&��R��Tg���-v��2��ˣ�b`�+��u���;w�׆]K;=�й�'O���8�{n���kb��$����AS�bc ���JYC�#�s�W����hX�G?���ޏ(Cq�0Ó�)Р/�+h.�<�ã�S�Y>��z--/�,,.��>�`\igr=sq������vۥ�yo��_[�g��EW�)�ґ�� v�ң��/lE�6b�_8q�Ćrn����xQ�[�_�\Ֆ1t��[j�W������+8�g�1�]�Y��=��wς����+�ցf+���{G[�;�ߣ�9:��N�sR^�h3ڀ,��õ�ps2�S�(8���Dy���o.��r��9�α��)k�����>禛�_��/_HZz��jji�;�pf�-G��@�wy��g��e��^�c:vH�IPxWy��Jw�q�ɳ��`!�4��?H�n���{��f9�ڿd���;�>���{j��e��� ������{X�~��k�Et����q���I�g��w~�����8�:q��x�-�^�|ߪ�Ws6"a)�w��~"��f��۳���x�୕��}-��ג���jjvs�Ѓo��#�V?����Ǫ.f��
=F.�G�� ig��w�AX���h?��};���},��?ӎo���_zϸ�)<������I˕���i��=Z[�ý�G���u�������z:�2�����8åA>	�E�Ҏq?� Γ�.�������K�F�'�u���x6y��������b�.m'��Nb�3�9$Q�EFx-�E9�4�T���B�t��8>ކo��x��m$z*\N_���_�)��=t�/�*0�g7t"g<�V���C�<������l!j�?-�������$|�{`����ɼ�㹜������1	�2yx>�L�}	Gnr0Xt�c�X�g:���l��o���%S���}����0�{�~9k1�Ɖ�|���I:�33d<�8�qK�7���C��e�K�ȗs��@�<�����oO�s@�\G�h�ؖS%�<�[E�!MhYf��H:�4�1#,�#�tC�_�c_��Ky�Ș�s~��d����Ȝ���pX`9�nK9�1�<�^���[ɹ,��a�����8�O���t%�j�n��7i�.s6ctn�l� �F��j�o�S���w�����ߘ�7&���#���>xVz!��t�H�Rι��磷N�^O$템��F������p�@�w�X���gΜ�?���q�M�\n���̫/�
.̞;��4�vf����h6�o�|������k�# �<Г�5H���A�r�����W��U%�BiӍ8@�!�a|6u��#G>�|W�.�9��Z����	���'��n��}�ǎ�����ѥ ���z^�����6�,�Y��ܘI]���G�N݆�[�x�!P�C��o���\�3+C������~�n�Х��r��Z�?��T�ywp	H����p��ܤ�*�es�Ŝ��O���ʑ`�~���f�!ǧ1�Z��Vi_<(�S��䛏��A���8��;ۦO�K������84;��~��pa���:Z_]���yC���mfS���ÝZ�=f���:?ڻgO������K�P��
ti�8]�m�v�؎��^{� u�9/��Z�r߽����ʹ�vxL�F᫼��m&2� �ci��W�/�6��~�a�y����)fa�س��N�>��=�����g=5qzcs�S��;��;n�����3&�)La
S���X�A�W��	������;����$~y���ӕ��9O���&ϗ��t�&���<]�'�P7�I<Y�=����v}�o|�g��y�q����$M�?��� �����)m�8C�\����,�r<�+��?�+�{ ��/��i�>��`agwg����f�����G�7�ƀ>��j�(Ǟ8�a�iX8?;��v�(��,��F�V|e����L7ǐӾ��
�Y[��B�'��;��L<t%��Hf�/�C�ø�{�4��{�q%�YQ>��w>������<�XAq$��1��k�g��3���ò��=G�x�q��ٍ��p
�������];Mmnm�C���8@�q�v����-XaR�G��@|���ǹ[�vg66��9gm9����.Ɓ�ŉ͔q.��;�˻á�������8i{Bש=��>���6�ɻ�0�������ٻ砕�Y][n��g�ӧN����5f���-\u����ՍճgϜ�?z�=+��_����[�י��:ڃFSx�@)�)La
S���0�)�� �v�*6}3��OL:feh�.�j�+N�g�s"�$�O�]�����u��(z��n��4��c9��7�1������T��p�Ze�Y@��HA��F!`fVޑe���.\{2�v��vj�Z��$9���:!97gB���h�5���3�x�̅x試�93�f�?�:La
S���0�)La
S���0�)La
S���0�)La
Sx&�`� ��2_��^    IEND�B`�PK   $�4W�'TO/ �. /   images/7789289e-5858-4b68-a160-e98940e09304.png (@׿�PNG

   IHDR  L  �   �Y��   	pHYs  �  ��o�d   IDATx^�`d�Y6�jzQ/�����f���$q'NR  �||�(!$�ҋ�`'�N���]���^$�z��G��s�4�FҌ4Ү�=����;��{�{��=o�\hF`�#���������Z��y�,_��[�~JQQ�8��Xg�a����q�^�H���N��o�os]�F��!6��L��x�)<�±����5��"�S���+i�5�� ~z�v;�g���`���Y,��x\ֳ���a��Tm����5�7�{N�������_>�G������ǎ���2X�C���(����|����ևY�K� ����FWI��7o���A��ꢢA�G+ˈ��� )%������֖��W�8��x]�ꊏ�U{:6,-O�چ���֒��W���s1��s?l�~��v�Μ����#0������	�~h���� ��J�����"X�s��(T�u�/�-y��ع�i�Z��۶54��3�>����T������g^�h����r"�j�w܅��0F��\�7�hC�᳋�ҒL��f��ro��E��\����5�x��^PL7���] Lo��:�:�O?>���w6~�>�������0F����P�'��x>*��1.�)�-�:w�\X���+�wlZV�{���������Ν;��>Tb^��c$Ϳ����ӗ^zi,�`�۷/���5�F0�ƍ��V���v���}O�����S�C���1Z4�rc�:��0�~�g����~}.��8X4�����y������G�W�.�a�+�ߊ�?O�T���sm��څ8�#`��R���6X�*���+��|���_�[Z�ڥk�t~޶�u�O{����9p���G	^�n %�l-A�qc�����M�`����Lf1�N�U�$R�T��p<�'�������w2��-�>��|m���O!�/�w҇��A��^�H��/�� �QlHY�7�_Ҵ\!h�'�i�rZ��*KH�7@��gB:K��#�����$�Q�{G|��S/P��,r��'�o�]��-�Cc����~�vb�p?u_��qKB�]q�حґpK[}6Ɛpt��^ϸ�A��td��%����MZ�Ḽ��㉯�6x�\���J(�˜!q�$��IS�k�QǟX��{�(�j���d�$�����?�Y	��5��B�͝n&�i�B�u�8��A,/vٸ��߮��ᡫ7����>�y�l��Y{��o��k�������՟�󕈙�>����C�/X���K.�������y����������	,p�|�:L��<̷֔�da�rӢ�[L�eLߵJO�cV� z�8�JQNS���FQ[��C�Qg	H�5*�enq��b�Ki�E�~Hi����q�r�o��J|� ���y_�� XCֳ�YbR/�RS�*��Ħ|�T�]VI&bґ�Jc�Y�1N���ؼ��GP��X��J�=*UEA�zK��$�k�1�>�̃�;���2�9����5�F�%��t����>q$�:,�g\�� ��O9�J$�ޢJ�H{%���V��;-� F	B_�������Dʱ��[�i��!�D��3U$��Y%<hS�i�^��.Jʊ�A��c����>2B��5��d2)�ᰜNUcU �kv6��9g�[ƴ̖���P:�6(rI�%�u���		:�P�.�T��.q���x�����;<%���i���̯+}�3�^��l�!����~ɥ/���o�) ��`�)�}�SO����������w�s����`>�8���ϟ�Iko�^��I���:%ʵ���p�J�K������x� ���������2"q��>�4F���=�3��N���UN�8�F*�0P���pb�a�u.ymGDR1f��#!��HKw�XN�\t�θ �a쪜iY��e���a�"X+��:��5i *i�� �IK�L^�Т3�͎��p^R�U�1�9:�H�;� ��H?����`���/a0�y��s���]��'�e^�x`IL�1F�2]r�+-_��Ļ�@=��+�ŇD�:��Ź_Y��ŖN�A@2�/��EVZ?�ӕ�[�� T] ��6_T�E+�+醲2�q��
 ���%���:�1KĵK{tS(�7ewH��#���=9�3�(�b��ڲ�l.��2��ƞ�L��;�MzC		���d�Z��U�B0��>�cp>�?��B�a+�]6�����[T������~��p�����΋f� ���5_��W�	����;q��M��填\���h���Pip$d�3( Z��h�K�d*�<��*!�qx_q�SQ�؝E�r:)G��e�@�#.��e8x��c&���ZOD���%�Vh�V�z�G\��ƶ-)�H�\�o�x\d��@SB�`qH��M1X7�����t�pGe����m�%뼲d�]	�l�Q���ф�8�G4&sR�ϡ,#��T�ƃ��MY@�81�8�˫m��2�x��G��O(�r�儴4�e[*,gaql�y$���9��"Y��r ���}�r�,]�̓?��1�SJ���"�`���H�D��@�x�OݴոӲ��j�K�$ ��)�L����8�E�NI��Z$
�]�n���p��X��=iY�	�:g��*�֨5�WΊ�y����6&őH�v/�@�-]��3-�31��V�A���y���w�,߀yOh���({R �^����Rq�8��R��c�
X��n30��ߙ������Sՙ��?���V�<�����V������;��%�0������߯@QQ��������� M�����~o����t"`/��#�q��m]��ƫ�݋�������=|��� fX>���!��Iw[R�����C��<���FiQ\6�Fe����r�K��" ���
���8��N�˱�1��NIxs_K8�]L�j|-2K]Q��<$���U����)���D�}��R����:��$X�_���y�V`4BKG	��J|���H�v���*K�T��D�-�cgkJN�I��$���9������3�giiJV�b�q�S�]�T�`�55�x�L'0��Gcr�9-�p!{$k^�O5��$��\I�w'eN�M��쁲+-1\�YT*���hǣ��䘿H�`�L:
�<+a�_�I�2oT� �V: ���h܆�9�-)�kMʙ�a9.���*�q�Z�l	������+M@�&�.rJi��든)�1�!�`���ưtı����k���4G@�[̏�e?}���/�_Z����杳�����	:���`�w@X ������Z�/���=;��ZbV�� ��G���PwBô��H�5Ynd~f~�b��n	��u�`\���џ��a��nȭ7�]�]g�,!n�R���
X�n�ʜ�B�O�_��ўA�%�D�[f��3q9�jT�m1���µT�,5�Q`�5%	�����^�r�[Њ)�	�r�]�����v��v%��|����|EҜ���9��� /b�����<X�.��+s�í���Wz�&j�V�[����>&���`/ h�nUqB�:�R����[��rlSZ>�p�'�'��z�e.Y��!Χ�R�
kN_J��+`�)L08��2����	)� �{�KaO����DEc�~��?�ߜy6���9s�.�=Q�$���MgB�� �s�1�[K�R�~�.���\��ι�+n��,R{�n�M��ڞ���8Ly��]���0+�o}iR6���ȥ7�a�r`/�}?���Xq��·���#M�lrj���r:rW���C3f���{s|�c�,�x<����M�bw��?��+��[���X�su}�����9��f}�'�Q<����X"�:�AϚB��8o�S�݄���BstS�&����a�.�(�[9�&���>0��Z"�˘֨�z4��+%"������V���P�O�ˑ����v�P#uy��a��)�XK<)����q$e>�k��r�G6]'Ƅ�l��=�$�r<K+R�-�M�pZ�C@�tM ��,��
���Ko�J�<X��s���%8���H���)�`A����XO�q躥�i��;�7㹺1+��Yu�K6,���6G��&�$ޭ���M%��啒�����Bl��ܝ*K��Me>Y��X���e6E���랛�5�=��S9�

�(,=�͈�j	J7�����if���ʰ�8���!K�;��mߏ;�X�IZ�pB]q+ܛ��	��*$Ow"�>M����wci\6c�W_�5�q�`-�T�We�<�t�*�"�x!�= KxJ�$+f·8��S}[Y���k���Ʃ��|��w�j���|�\M�٧B=k�e_��q�7u]����rR<���Pq!k/BFV[�д�Re� �dy}��?*^ �#����J���#����U���&�,��,*�} v��$[�8K�2��@�-܇�	��P?�� t�=�3JYy��D̓��3a\Ĵpn�pRf��v  �}�:� ,dā��wi�x���Q�C��9�H Rcj���Q��C�m���}Ty`:q�/�4�¡	k�|f�� ��И��s�zU��ua̽���r�&ݎ����xA��%��V��dS��"Y��.��`�|1jL�7�S�Q\�qd|��>;��`I�4,F0}�M"���i$�;+����r�J�2Nf$X2�!��P?�7�S������"N]�@WِH),UH����j��e�6���#-J���5�T��O��f��Vc^���K`^�)�2�ƕh��\Ue	.�5[�X_#c����zT��m�S����l
���E��wIEy�,A҈�I�����X���`��<~�ǻ�U����-L�8)�f3���{�9��|�ϟ]��ܢ��$��y��/G�����ȅ���!���/�=���8�,/�:,��!%���Ka����歲}�F������R��|�SB���R��""Ou{�n���}c)�u\��`��&2�2fIϝȞ׎�}?~ZN�<#�M=������d����^/��w�5�Cg���_��Ψ\��K��T�a��J<�.0�T"Ͻ��X�\��c�a^ca��^�<��n�����tv����%����~����p% 2ښ� ���Jp )a�kUP�_�gV�d3��s�@���
�D��z��3,K<��x���O~���<ݨ�>��"����\$�6/�u�b-��:4�Ij�q�m.9�;"+D�<��mu��,-N!� �S�ceU��Ί9n9�)O<�<��s�G�t��l޴Z����e�E���\7�e�y��w$AE�0Jjj�.G�ᆲ��]H�\1�R�!�tҁ��z����������Edn]�,]�P�{�\~�Z�a�H$B.^�u$�#��eCV(���I��5(�Z+�-e1P��d�ztvĝ��Aꀄ>tF~�����+$D���a��x�Vy�;/�ʪRĮh`ʭ_^m�;?�W��H<��V��榲�� ��Jl(�aO�e7¥���O������#O>�G�:"~��#s�V˶m���6@NUc���5�� u�V�
!5J�T ���{!\�S����fC�ȕ?x�����gG��3��zq6�����G`?U�9ka�g���탑X�թ'���ڃH�MHM�GF���Q[�Y��/�P����ԁ�VI�A!y���iy�W���J��>	�T�@��1Wm�ɎǂR�C=�YG�n�����֊�nD��q���b-���zQ����#�{�E�OI�<�o���������r�=��]i�����N�3A����=����R�W�jw\Z����.����0[�}ս8~Vimj�������~�ST�pB-'����.�<�S>����J1���8�ň�ٰ�-��T_�N�وE:�SV�����=�`9Շ	�DR:��~������@:�|JS'�`pgSS�<���3�r��_}�òb�"�ϣ�C����{dQ�O��y6�H�%) 
����nEv�l&�W�����G�����ʫ��PV{��G_�x�<��.Y��A~���;��fd~i&��j��]h��}!iK���Ƨ�F���j�@u��sÝ�X }�2DBH���/��}�>��`�ϟm�_:"��ޯ�7?z�\u�Fy�]W)���@f]-\g�oC��#q�<� '�S������Z�.�E��b\ͦJc %���w�c� �=��tt(��1%(���i(P���'w�_��ob���M*���bFۙ �rB��4���o��W.���LMZ��:-���o�I(H=ݴ�����2
�����\q�Z����%���L�~�U͵�ꋱ��_��$J��/��ʻ�ݾs�T��o������?z�ʿٶ�Z�̵�,`��l��0经����_�mg`��j)�N�[6]	6�!+�&���^y��I��-�UIwX�Ah�!q�RZ�@L0���YZ���?Z���4��$L��r��*e��!E���?�e �k@v���T���V�!���ny���ċ�ōC� ��ۍ�\1��X\��j����W���L����HD�l �h��B±E��|�&����^�"�s�Yz�g$����ny���Ap`n�G�(� S+-x��8��/���`I)�/~�C�� �r�M���ʙ�1�<����|5x��rWP�Y��� Kt�� ֤�GO�C�=.}�~h�pw�S����$�9O"�<����������ZU5di��o��#���mqiC�m>�p���E1dÕ��2,��ѷ=/�*�>��8pB<��X�.�����*���/-���<�Kq�Wnȋ�bj~`Г�oż����3�A�~`�s�c���\܀�*fKc-���N��Ϟ��v bv�;��p$�ֳk�C���'��{
��G>���>Z!`��|����6;�^sy�>�� �cj�Պ��X?�8n���/��W���N��K�P��P�?
���/va��r���r{3d8�K��VmrJߎ ����� (���ҥ)��@���5�aV�Z<v���'�$�4b/q�'%���b���/�?���������;���Zm%]�ݭn���)�xfoQI�`�0���}z<�lJ�5���w�/��K�f�߲����|`�m�5��4n1�_����+EM���<d锩e��A���>!�>�l^� Q�Y�K�`�-�-[��ŵY�� 
����[v�|I^�������v�*q{�J�sA8���Bv�CN@P�듻�gj>���Z(ؑ�n���ޠ����D7xeAC��c��z䆛n��k6Hee��`M��}�5�g���������n�#�3��nX�ܰ�9���ܭ�9˔�E�S�%H�_��� �Y�٧w�s��)�`��T��|������"\(�s��}����<.������O�7����r�v����ʕ�ƌ���=�N��㐋 ��[���Wps1vŴ�����+?��/`m;�yt��M��ʫ��BLp]���vy����ԩS�x�Q~���O�g��^ܙ=�Z<�a��H�Y}�'�wpR㧰u(�SK������s����/�����n�+(*��b���r��i���k�ꫯ�%���^�����X�P�ͣ54��B���m��[��In�<(߈d��������˼�~W+��~Xd��m��ͷ�KP��Ϋ�eWW�:tHv�zY::�Ժ&���O6oY)�^�	�N�=y��;dUw�7�,ܦy�'�-�D��&�-X� ���F+Qks���g;d�E��o||=@E)>�`|�����r��qXA�0fI��<��k�����pq��p��C`�@��P7�}�`����'H��J��aX���T���^Mh>��q���w�G~c�zn�@��=یq܍5٤�\�B�בC��W�=�q��3�y���t�Sah:���U��m�F��u����߿<t�_�Ͼ����n|z&��LX�����������c���~���w7�^U�;��p�|m
J#���Aٵ������))/����`ť�O~V�,]>b�n���������C�E�PP����4Y�~�߉�1^,��T��<����"m-} !��6@	�z����t�b~+�S��Y��7oăn�����39u�5y}�>Y�~�r'�lcL0����e>���t%�w�+����Pg�V�>؈������q��o�O~�d��c���C�-����Ikg�ߨ�r���pKy��4/��|W���
��0U���J�U�+�nk����"�Z��������c����|>�D,����]��H4�E�;�� ���VZ�@+��ݱx_5|���Ҏ}R��-.�[��������#_�����?q �CY�z�����#��3U���s��� f�����/�5�bb0�Ups-.O =߫��P, n�|#sn��������|�ga�0=����3p7u��������-Fi�+%�]^{9���c�O�Wh7�~J�| �𐢟ͧ:%�Z����˖�.��	�hO>�<��C���s	w�)7ݡQ��W^9�⚆�@9&$������| ��J��&%A�m�����A.5�[%��໥��z����I�����J�L�*ʉD�v�D�F�*v��t8�u��޼蘝{��� �n��Kw�i��7~q�����M(h{���4��,����ӝ��N4�N��1����%���*��u��B�yp��Mp�L��"�.�r�e�Ȝ�Ur���ں�cnH���9���_�lӂ�ծ�P-�>���ލ��`�����5%<�ڡ����N.A�r�����;W��_
8��NeU��˿}Y~�oIc�>�����jK+s�:t�ΔD�PR��&u��b�=�୛LI9v��=�,5U��w�G���RSS�u@V�\%��������'O>��|åRW�>ċd�Jmqy�Q�/Q�.�7�=saA[��'����pSuq� �vE���}�+_�.Xa*ծġ�m��,�$���g���pա8�� ^� (�"�q�3����ԋ��Kc?
�<V�VY�|���wY���O��{��[��{.��[G�u!:�����5��=&=���n9x��\�m-. ��n|^j�-�D�0k��qZpT��a��V��'�|����k(�.�r��Y�N����V����P�N=��^y�{o`Ԗ`�'���|��p����ɤ&���X�n����HEE���B��z����\ w���� G �[1���_:@��
(JH�m,���}N��a��4+�W����W����a�Ee?&Kt~�r�f���������K�駟�'}����W|	ǎ5��8_Ֆ3-�,�i��Ҽp�4G�t6�,|dg�������E��y�_?_�0�x��U[���p�Xa���*�S�~�/�du[O��$t˹A@�Ps���&�2��	�(����D9�J0Y*������#�kX8"��|���b�C�^:��n�.��aiޗ�X9�����2G}��!��ӧZ��g�<���&˖��Ø�����1��m��O@�Bi�l#�40�����ZV� ]p<��������6 m]�[w����?D,EC�>�N���/�����H�����<�����4�Ί��~�B܊iڙs�@-��w��k���?�r�M�bNK��|A����z�|�K��^�?IZ-Kᖙ���~�wo�\Ne���9��Yn��}r�{�X.��ux�n/�������o|��"��ҫ-��l���l+;-F�y9/�[0�[�����GV��*%��⸍n�]uu��������� ,�@%�b;ܣL��2@�2�,���JY�F�4�?���U}]C���z�]w�?b��6�c]�ar�ki�8gt���p�zt��v�I(KVd�I���A<�ݓFuQ���uAp�������7�-���N�X�%�����.X�{ǀ�K�>f��7��l���9¬V0����������y���|���r}qc��+�iT����|$����-!(�2�_F� eԦ���E�6သ<�%�`o|g�t�`fV[����X�=[S�Q��w��`'k���=;��k�� ����@]��㨡�-�JE��n2N7�ͯE??pQ��P̝[+����e���Faь�M��C�.��p������?,�m� 2���w�y2%ߣ�>�8��u������"����F��;�e|�č@��v��$�6nV���-��T>Σ1�f�/8�tkUW�!XVV.��������߫���J
}�Ӣ� ��(ۤ*P�C���;��'��q�gׇ�@���XB�������Yee������Z���ý���s�3k��C�9�օK�;�O$_��G���]�#�<�1loe�4�a)�WMiTx�^�����i���7e1�L�lp��J��OwKBř��S��u,��uk���!Z�|6ÃIPV\f�5{G��r�)>�����D����*Y�bu.�T���	���N��(�C^{�%�:Z���z�)���d9�z�����O^8A��d�EI�rf+�ls�Ǖ��@O�	������@�x�sn�]s�u ��S����t:fZ�6�,��إ��\�.ٺ�y�:��v&6�BAi����jw�X�@��p��ɭ�X��{`�+A�?��FrN�v�����lـC���7�Z��2h}��BwFS��ᖟJ��ڡd�!G1ʙ\ښ5kd���:m�l�g+ܔ�{`�k�s�ąk&f��"���=��}A!����WKNn�V!fw�8��<C�J�B�N��2(/?A���#b�@q�pU�l�Ukr����Q�7�Ș�)E@m��� @wVL����*���h��x�� �8sod��A��]�)")�\̣��Cy��
�hG ����t�mڴ�E׃� ?c�q5�%ZCf���C���f�S��'���6!XQz��I��ƴ%=j1�y�5k�ʆ������xP,���^R'��3�~��g\_oLB���mp#��)�A�O#G�֭��Sa��V�eg�*��#˻D�R1 8)62�\Z``q�Z˵����fN�,���H�7�O/�#S?ڵKdl�X,0��6Y�54(�6g���䛌������F_,�4��I�9�=3?�;$<ڌ�O�����ɕ�b"����/c���Ȳ-NJ��I?�|�>����9��D��o|�ߛe��zC�?�ҙ��y�;7s���VL���g}Q���c�����:U�6��Z���)��n�C��Z���.�����n�س�~p�5�3�zO��6.�5��g��0�Na�!g�)��Hɾ袕���\�m3 ^}N�����KN�F�?!_J�AM����S��1 �-�B�Ǵ����6���w� �ܵi�L"٫,s���|4"{_
�Y����a���9�}`?k
��0U�l�s4�px �;�K++�8����M���>��(~w"hW�6v�d	gb��D�T̤m0�Xw��S�� �~��y��8���2��<Їa%��ѕ����N�m�[��ċt`�r���/�[�v��q�6�d�Z�/%�i\��Z律t�`x�\��_����� �M�s�Ҳ2d��d��߱��a��l��'��Y$��Rx�r�wc�˩�]|�W^ꔰ���ra�A��5i?׶d���Ƥ�;�y%(Q�*s�%b �B7B�I;p�/��|��L-!������b���B��~ |:���/x�������3��b�y��j�����Bs� Y�t���v�B���IH9�����j8Wu���������>t����6�b��)�z;R�M�&�q���&w�s�<،t�,9�?!�n��A���a$޴�����!�N�XU	��&kt�q���� �V*֓bl�ō�V��`S�3��`d%0��3��h!��3:ikL"�<-} !*�!���&�l��/؟�5�A�]���D�R-�sP�?�0�]������o����D���iԥ���*Bߞ��}]�',7H/����^ Ԛ�n�Ný�8��C�`�;X���������γD����PoG�T�����`�M�:<{r1I � ��d�V���{c	p�E0�t1�snh��G� �O��h����92��c�N�b<;`� �'��Mr�y����-��S��(~GΤ�{c(j��(�φG;�y"p�e�%���~��ǒb5�;��X��~���5�|y�4�;��{�W�%�q�:�qR��|�U�2t[-�4eDh�Y��.if7!�`�
N0�3�zA����P�R�a$�U2
��9��޴�d�ɒ�ǝsż��K'Ò��K�%.��3b��`���Ir�6�❋26(BA{�$�Uɡ�$<�ieM�"�y�|�}���#��
w�˩�urI0�;��}����^� v{� (T�%W*E�:c������P��������<_����t���Y3Gr�ZA.�D�;���.��>t�䩃�b��R�b�!�����=�o���h��@�^�v-�nߞ�ݾ�[�����)4N������8*�_�J��0Kkg?5����g�X� ���D�t��Q|N�>�O,kw��"���0�kb�/ݨ�BN`��8����#�d�ĞGey�v0e�����4l�z o�X����E5��L��P�<
`�3���K�ވ���g"`&p�,�/�ʪ���Hӱ��1�[�C1�FY��\ �s�bZV H�)�/[㘦1���u��O@بOGe��-m84myj�N�L-���׃��K�P6���o<N��x�9�����x� ��,�{�] ��+�{����5�C�`$����S�����(���(cL@�����`9�x��5b\��~�৉�xL�aklM���Q�ҟ����? ����9 �^��U�~��I�i?�t�Y>f����N$X�$ �^��Xs��H��t���%U,��Gn�|��98��N��[Q�"��{���ǈ�c�=V	Q�ZI��?�����*��}�=}�����8����)��1 �ț���{�9��W[��oh;��-�3)��B��wu6���y߽7�����g]��	��\�.�(p]�k[����7��~I��)tX��A��`4 IL�IKe$J� ��\6
�U�w���V��j-��#/��U�7s���#������<������T�z� ӏ~����9}�l�E踛�	���@A+���)s��ϔ,0���ded���Y��Z��9����@�0�  ��w �-��%�xj� )�ݲ�� Pzۗ���W�Z�o7�|��L�x�y����c+�����+��ʡ��e���.��m�H�P\�|�t�9����3�<�)���^�S���2�bt��F��'�BG5ZJp�Mfe���hHs�u��f`�~k� #���0oEp-���4��8��"X�
�$�O/���#)�d\@���#�M���3�B�6 CX��ZA��.��
�n�E,{�O,ڇ.�A�h��A�ӓ�"�ۙ��X/�Â��6��8D%&'0��{�����bHt}5=�Q��i��Q\���ȧ�&bA`3��74�jL�Ov�s�Kx�h��R��R�P�هIpY5���+�4yyp��S��Z���+��-�FlN��fN�(Tɝh,�p��뙇�x�#� ĸ�����1?��C�/�IϧU$�>�Ƴ�F#$a���5% ȌS�U���kKJ�\Yq�7�+�cv����;6�.>���ԓ�\��S�^jſPr��d�F�s L�a���0g�k����lB�!6	M�z�5]>	@�ڋ����N��_+�PA9V$hx��Kh��$�\���ɢ�K�j}���(^0�� Z�������~c�B��5I��T��`z��|e�T����F�!e����;-�)���RҰ6�ve�����TTT�����8�zzI=(��l���<o���;^X���SW?�b-����m7~�oSuQm�d6�'bAz=����X�xh��&ӅR-u�(�zr��M����ַ���)���	^���.��}����ʡ;S� �wG�KðD��
U��!���(N�"K)e�@[C����t<����(6�H��	��j��<��*Z͑.֟s�DG4�c
���E�Z),�8��JMC�,^�b��u�7ݠ�Z���N ��FWS5ڸXl!��yh���E�t�8���[�)=i���♢����qh��_����ٍ*땨��
2�U�Η����P�ZI?��a>�\���cEm/�m7��P�oj�]}�A�G.)�#$�����_��s��|F`�hRu�R8Xcj�X1��c ���AC�4�6@��WiKe'���hb��a�_$��4�7u�����?�R#v��1���*"72��}eڼc��d�Y�X\2�¨�0չW.Y�[x��:|�_���5��'�f�Ö�$�x�Eq%�L� �6���S3�O�  A��;p���&��O�-遅��8������t{�=����& �Ԑ��݊u��P`�r�H CV�L�SPj����������_n�z��Lt�q�1��5J%�c�+�	\t5�D��X�xGT.۶�|t��\��� �������R������A��A��%��m���W�UT,;�Qkô2���x��E~��2�wUp�ր����fbX���-p�G	�Zw�VY�g�$JQ� �W?�D�������������ӑ��>+��w�̩�8נ��<��]Z��^�<�ܳ7������7������'���>���}���7������n��P�+����M��zNM�)#r��
�T��2d��si)�Fǟis8�������� J��,��%;P؍K�z�� ?[�U�6�K1 ���OF�e�;,�{�(�kE<@�Qh�ę�r%��"@���!��ҍ�BE�p�?�s�9$��}�+��:E$�;�a���㑹�t���e	���*4K7�eb6�vఌ�U��0 >�
CVt?�15��sQ��#'O�X,0&����8���ﰖ�	�(���*����06PN݈�vAn�W�3b��Xq��N�;���%����4�?�l��9�}�}�`{�_.��:pgX�\V�#��x�r_�����Z��1��8��?E�9�z|� E���rrO@t:Q�.#�o*�ʻ�\K�݉SA�t?��e�����EajXF�K�&0�#I�L�����K�Z=�z@�B�9��	 |P�Hm���x�S!���&��dD��RU��Xu���c_����yX��*��`�:���ۇXȎƄ;��?�2��
ĭ��oFM�`�o=���� �żc���ń
I�fbH@]~O�������Z�řV.��*T ��&/vx��>5���,��~G�Z68���
��us.�;o���_v�vH߱m�ϸ��;�Q�rū�캥��ɛp�U�z1y�c��I�����Y��Zl�QR\�פd%L������?�������_���ڬ&,0�Ν/�w,l>�~{_�(��\� w��u��n��?���}�K_��TG�ɗ�����^�8��
�(�J����[<�Ťm���]9_ŵ�́yx�F��<��ç��z��20�����֫�W \!̜�*���Å�,�iJ�`�(Ф�28�� �LԷ&��_ <ʲU� ���T��/���A ������S���fh4%`��5�<r)�	Ծ�!��1�Ҩ zz��;m�2|Տq��(�[�8�f�e=(R�EO�'�3�+&� ^Ll�W§���ܧ�?ٗ!��m��` �����e
4�zh��
s�8TF�_�C���.�JN`*m8��UZ.���w:d�������lc_��t[���õ�-�< @��0m7ǉ�TYl`�=���cr��|fE���4������m���h����Ul����{����q�}Պ�����&���>9sA�>��x<�Z�YK�@�&�J�u��G�d�Z�v#s5��;���B�&�I� ��*���	�7Н�����v6����SԚ�b?�r��ge���3A�>���.����C���>���L�� �cp��@%��{�B������n�t�9�T����8��K)�<N{��[����?ɡCۯ��a&�����?��w����~�������.Ќ�[V����O,*�%wB��Ҕ��,�^���L�����`�_~������=�덦��s}���Й���h��3�^��e[V�Y��B�����o~S��K_B9���v�5����������I&F֙ADXt������JY<�t���=�K�I�ϥ�6l�Meq�C��c0$�7zP:�L�*aVg������	��Ҋ`�S S|G�C�<�bZ����t�9�4QF$5�H(����s�N���A����+&�ܲH��J<�������ڋ=8,�8p�2\0G�[%�=,��G�x��L��8#Q�/,+�"���9p+5��uD��x}Հ��d@�xчu���V9[(O��A ���"�X���7��	 �ܬ��e�iY���OO1\�Ŵx�l}� $z�O�H�R�[䂕�X~���k���Փď��i���#��l[E@�T���	���UR7������"D�g@�Ј�~XW����=��œ�v�,�5v.�y����0���pǢ��gciQ�C�	'�����Ay#X)�Qd�N�e8��J�P{	i [*}��6.+/*�9u�Q
�8�ƽb� a�1[��&�p�C)
M(``���*�+����m��t%�~���Je���$�/�g��o�%�Ȝ����.y�����~RY�ȝ�::�њI�{�Yv�g޻���>������'�/>�>��T�Ӑe.%e��-ֺ��C��4�q���{:���M�_�ܜ�9
cN����S��>��w;��m��-�}���B-�|��u�ڤ�+a���3�nJ�����Cn����Qh��gs����neE��|Pڐ�F������#^7���"�
��ɣmr��qzU��+��p���t����8P��qM�vh�	.�# ��	�6,Gm�$�j^{�'�/�Ȫ��:m���g�u����/%H��B\�.�Az�O�%6�Ն�s�je2�q��25Z/2��o�~6"W�21W|�h�C�ZK���݅��^q�P8�a��p�Y�Q�W���D�h���Rv��8��2LȒB�ѿ�[��h5i �~̌�!�Ζ~@��ׅ��WSe`�eZ8�9��Z�L2�h�=e?����C�$,��p�����ę���Ol��C.�
��D��x�''����EuO/@��X�ә��K�S��0���*.'b�A�˺KK���DS�d�"�#X�������[V�tO��d�T����k��0���0V(�:{���B,b���EC\Uc�')ϰ��`I>�.72��r0�Az>��0��<9(C`�k
{�<���8b��r��5R+--�CnJ�:3z���&� �8� ��xK@|���:�
�*M�.x���� �r�Z��\����qj|�#;��}��X�N���J��&�*�⍷!1�E���
��Ƿ�8�ۆ޼��+�8`:�X���O�7Z?�=qGQ������$���[�R7ӑn���T�hxN(��G���6��B�F��N ��h �0V!���
��w���A_,uK����B`kgkX�`�!>9�,�[�T�"x��dp�"� ��r�A &7�xG��=N7\fF x��@��kYV�t0!�^��id]��B��t���A_ ~�3���M�������r2`W���E�QY��i	��;�ax*�R=�!�N�h#S/2�v�Օ��W e�:H�;�_�L#_��I�ʉ7�!�iľ�	Z/P����Բh�A�����;s��5X�v����Ųb휡l�����T�|?,Ia���QЅ6d-Z�������tQXĦ���� �e[�*�vW�%�;�A���tV�.Y��Bj��܏����X���owSZ� �<�X�f�f����VcA�p<\��:�3=�W!K`a^���t���~�W�cl��7�,<��I)T��L�>ܐnyu����~��m��50	����Z#���I�;e��r���oPak<�����V�X�B��~� ���'_����6Ȧ2{R6�}�ʯ}�_�[A l��N�"�kɩ�{ĩ} H���H7���h�t�J�T���H�����|���s�+P����yy�g��X3=s��>���<����?�������h�IB[����$�����{-��b�&�Л�=r��	���?��sL���\����s��nߩ������g;�S V�^A�X_�/��Wɜ�������o�3]r1fj)�b�鉐�_�NY��]ؘ(Z���C���d_
7������ ��͎�.�Ƥ�S�e�"��%�:�tA�1h�'B^�!��5�qV-	���e9�5�W�6�3<[Ӏ��q�T �{�'"	�����K�qĿ�`�������A,ֺ��PS���������˘*��N�,�屬¥�V{#�6���2�$G����>���/�I&oC�G��-�R�Ct2�?Q ��&��|�_�V�kC���>��#�Xł���aU����IjP6�.sL���8�I<���(\�ӱ4���k����B?+T���b�?أ��m{�C*���ӈ�j�oJ�s���e��b�����u��h}S�H�����9U#�Z��z��=�g�;)����l�� �O�Jc����pi#�J����z?Y��Ҳ��ޮC׭�@q Q� ���jJy���מp�x(���9S�4��ϩU^d�YPz��������7qpk�	��N}�`���qK��%1gt����`)3�Ϡ(��t>[� ��y�UǊ�31����^��C�g��j3k�9p.�+.��@L�P�~�����LNv��0=��s�?�h�w;�B�՞ƪ���9{��d/����y s��}���� "`��j��a��e ֐�0�4���<Š�錟Ҹ��Q�BWW�Ʌ�R�C@�����u�&��I��1>� �3��n$'������`l�Ӥ�G5��� �v�b�{<���>����:��� <� 0� @���(鬮��-d����pMr��Mڃ��#�*�Lsa�܊e�$�0[-Ӧ�~u��8����e�f��L�q!I&�\`O'��81�i:�a:(�a �NX]8 OF��ۘv�cĮa<a3��`�2�����(�a�&R2��D�o ���Z������cxw�Q�+����Uʪ����͙��nI!��t�|�A>��Z	3ׅ��P���à�+Z�@��rD�& ���^�#�)>� ���c����έ1�d����d&Y�2;a�d+��믺�נj(AF������Z',��q�
�4!s�r ��\YT�b���g�H>�R�T� ���N�ةw�	�b`�7��C��`?	���j�<kt�^�ыVռ6S]������s�-_޿���[R\jĝB��ɮ$vV<� �@�1���<;�yq����O7�]��t��1�^L���v�W~v�'���2�1'�H2kE�<��mz9�y���t���+��nޤk��P�W����]�Z��{2�@Jp� �L�=ftd���ty���^	B��x�O��Ф tAX�N�B+-=�+��� bh��l&�"0����Ec�i�B�.dV������i����p*o>��T 
]� 0ʦ���,� �?�.���`��E )��L4���]�7�n����g�s6���C����>9�FkU���t��;j+��c�V0LX�RXC ���RJ!�6<`s�W}X���u�	q�C�@��@�h�)�x7u���D��j ����Z �i���.Ӻ���q�P�d�&(1�F�d���#pay`��Qɣ^͸:{b� *ha��Ne�3-Aj����-�m�K��Q�-Ѳ�����$�r��2oa�˦�M���N����ܼ�bF�܇�c_���m����ҥ��)\��n�OJ�l��ǎ����;�§�M4��v}��Y�`��������As6��;<�:���v��+���
����$cn�b.o�H��B���ÑB� G�N��Ihx�����FQ������`55Ӊný��e�?�͆Ö�����2�����:�Ԑ�c6����\�� ��O]�Jd�=��(Kܫ��������wRY2��죢8 eD3��w�&��T��[2�LיԖGwG�nU�UӢ��K�.��x`�|���R!
��cA�)F����&�M�\;�'ǒ�/�"-Xʡ��[��̆��D"�d�t���������}��[��Wr�@�-���ܯ @,/u���S���ǷiӖ�`���n�=@��p	L����?�oq��{¿�����'�~A%���8u�+�:>L��6s#`��e*7�Aڣ�M��$�L"� Jt��\�Η;�q�4�	R�96�Aj�$!p�c8�S��M��Q��y4/!a�e�&ZsxX���6��&1
�gf?9���MD3��s��k����$q ����E�,0�_�ӄ��c`Q14�2�Յ���+m���v}^�U��e����S.c�9���S��R2�b5�'��`駛4��I�m�5�%��s̴l�(h�b�2��L�=s,��MUIP�h�!ߍ���PQsB�̆�,���5��Ϋ.>���ӹ������K�=�`��a�S��$��	!3A���N�l��3'�|��*�K��������������XLg^����3�t�������FT� ���x�Fьu�Ao3�6��B��S���>s���@�3=��
ӄ��.���g�G��L�N�A2^Ԭ3]0l	�J��F,����ʥ�~���PL���+05�@���""<č�TWnA�Ƴ/ȣ���bT\J�IƅY�>�K~�����Nd�D4�4���˵����*�٘ᜬ{��Y>�a�0��@\ ���F�+�U���!&Y  ���8�ڎ(���^�i��0搞E֘9fv�-����g�1K�t��y{tU����bK̬�B<o���A2E����1�{���뮿��O�x����D��M��`�Μ�ߜ�橭+p��<zr�Go_���V���k�5�~��7�$,q�2���F����fC|L鬕{�Me����9$� �I�)H���4Yſ�Vj��|8N,�K������G�%�\s��t14q��dSE)��h]�0CM��� �3y���r\F!T�'� ��'�mf�x��,��H�ns�P�˚�VB��g
9�
܃�=K�p.9v�2(��G��e��:=-�q� �e����; �(�/��r�Mk�?���}:�`�2t]�UH1�r��i����ˁ�G� ��%r���@�e�rQ2~�bE6i�Z�Yi��Lh��<D����ں�*�r-�l@�*e��"���3���Nb_�@���
 ���E������J������~{VY�×����f�/{�K��>�f8s$���,�"W���q>�YQ��7�׿��Ղ ��v]{���Z��O��,�@`+����D�[|:��F�����:Z�&H���[ʾY�M0|L�g�Jcu{_2N�ǃ�@
�L[Ox�2nUs�p����{�=�M �о�'~�.!(  `f�� �8V1��/U���@��w���8�A`�1�X��N4��C�Tv�7�wnHK&gګ�O?�0L���~J���o�`46�VqW�A�W����$�/�;Lr+�<�(���yy��'����8�aeUߓ�7�� KB�D�����TF Z_����L��ե�	�����+�H�=�X3���
��g�9;�d�|)�E�sK˚J`�R��kx����j��4˛�J�lە�����V%?�f��0�h�Ȧ<���v�]��m���7Ս�� ����mg�A�J�T�ԥBZJ<�� f���*����������]]J����2�"3,��J�һ���=j�<�ب������_)�[r9�#��l�W��s��a�Yp�5syߙ�����&�̳L-��=α�fFZ����c��7�شv��~S9�r���8tZ��b���d��nZ.t��a�U��Y�iy�ݿ)��������e+C�7��U������!Et
giN�0�E�>H!�q��K��xYE����%x� ��繛Qbg>^��~���@��43Ԉ�ӊ@NK ��ʲc�b�q��vӠ	��K��g�)r��2�L ��ThJT�Az�
)�3�%�9�^o	h�;�_0AYdqy�Me�=W���é�������6`za_W��~��U�QKL�9\4�c�u��^�u_hS����ҥK���+�`M�I-�Fj1E�p���n�����J!9��V��K[ګ�L>8���a���fKB����ƹ�����6R$�ɲ�o����,K��4q��%���{�è�>�}�\�>�:@�ƅ��25�j����"l�vEaɊ�Ḃ��\����r�uH�I����9�3��ā��|e��)���������/-]΋e ��gU�(�CcF�A"擛n�A�.�,�==��3/�����]��rR�e�q��L7C�s�iWs�k�ܨTH���L�'�)/�0�p* `�dO�:��а�{��̠R3���ތ������r��-��W�+�J�#�b�u��e��_xqL7�ѡ��Eh���5#v��R��W�>�˾0��i�#���xCf��T��"��E�-@�TW�<��5�|���MA6o�|���#gΜA�Z��Tp�o���؃2��C��לҊJ⌇PC����R���S�M`nUsnV�xnTЧ
���;C �#��̮�<�=��AƗS&kf;ݑ��"iMӎ@�Y)�IЄ�W6�G�~�#5[M�]h� :@S��wN�
�k���+Q�:��;�NYA�w^���t�Y,`���)�C?��!�qP��3!ɽ����n��"�9ݮ�sE�}�����OJP+��!iTIr��R���"�޵�>���%jmP�c�����~���T ! (?��}��O������kBL��s�5��I!	�-�5g]C#ޒA���̸��O��%P����Rq�����\B!��;G�8�����-�Q/	��3���޲�����J\4�%eXK ���=;ٻqO=�{׫G{�y�*���L]}�Z�-Y�@�7Z3*}��FJ�0���~0M6k9|N�l�����X�-_0 ���̛�_�un���+e�B�Դ�W��L�a���k���L�ṣ/��{z��?�.'�7��e��IiIňKU������qy�`dD��)<v��eȰ� T
]Zrx�4�����}����B^�[�j�3M�G��S�i����� ��80x��ͦ���w֠))A�0��	Fp��`j##5H8g:h~��W0�?�B�cY�s����)`��?M���o�4�@�ة8�s�13���qAD�3D�d0
�k�'��p���9��ATS�������h�0o1�]t<�
�FgB q|�V���������Ov�|^N�:ď8+��!(�q������6��H^�5E����.7;�mh��@5�C�I+O:فY|����&ܚ���՚�%K7l�U�'[������*m��L3��gE�P���>��m�+Gz/������S"9X11g��1��:r�b���6r��z�jY�b���F�ܬoE�h�Mo�`��T��/�~R���+y�g��▯}�'����G�N �̒��4S�a,e|�z<��@P�u�F���wgo������3�D�<�2���� �c𦨂���K{��E�Hw������.]&�5� 5q�Z1|�z>񊥕q�tzƷ<2������6ŋs� (�
 s�D�[c��DЮ��1�tCQ�$�5ARa$�\�	 %3	����w�(i?�N6v߈�h�k�k͇Dk"��������b�C斗��G�\t�;�;P!�u*�6�+�k+� neY%��"Օ f����z�P-)�L�YE�a4^ØH;�E���4�K>��r|A�YІ�������$7���K��B9��>�Eٗ���{���}��g�L�x�v,j��D�`��jų99o�g1cn�r�ר�L�a�ޜ���y�e[����k�?��0��ny���{$����O�c�z�#�����\_�8m���U���+`����GS_���wu,�Ҝ� ��;���G��W°N̦ZA%˶p����7c��f�t/�B�Ƌ�pe�l�s.{z��9]�*.AI��q��i�iҧŉ�b���X&�tJ�����8�*&�X��hp��8�	Ju	#P<c+���8���p�EuQY��ˠM��{�G�3	�KaW�agX� �*X�x ��-�5��\��M��em(I��/H�3�T� ,��Jx��@�� v�BQ��=zD�2�7H�Z����u��XPQ��l���B]�HƫMS"���t�y�������Ծ��+��<�ma��2��Գ�L.<�\��FT���
8_;��˩�L��SpwuH2�'��尮@#V������3��ݧP(]AJWDΘ,�!fx��]�o�	���&���tB�8�!����l~��{�B�2^h��7�{Z���o��+�%�}d�qkp��W&kITY�@�z���8�52������@�pA�*>-�t�堙��}K����hE0-M<�y��@7������O
:4���k��o��9V*�A���� 牁�V���_��a�Lt��%MnI�"R`�36SI}P�C|�i����O'��W�g�@��Qŭ�~P�w��'Ǝ* l7���(Hł$��p-�����/,�z��/�-�H`�q�&ф"���
�	d�T\i �T���pN�b��Qȳ�Kߡ%�Ii�2Y|�ǥ�t	dZaS�X�'[���Ӎ��~ј�)u~�/9|������B&
�K��n],������c��]��WZ>�����|ڧ�v��iQ1j��D��j?��?-�������s�(j�F����ƃ,����^9ݝ��.d�D�����5��0|��|���*{^�/�Kok�V�`���b�Z����ظU�H�>q�M�|��馏�#��@�_���vV&��%��J��G$tv��M�FK�\���H���ҍ1eݯ�ŗJy�f��5�n͆Pf�	~�Ȯ����Z9�f=z(�|Ƙ'E�b�
7�㝸
���iv� ��# �(���3�3	:A#�	�.��?���И�m�4�fx�W�R9҇b�h�L���g_	�Nw���Yp���=I%TD�J&pRnjX٘XAn!�喽Gڲ��	����80��2�Q��@��Y0���s����)�������m���(P5�G;�k�b���a9��gr��O�	X�:䢍+$^�H| {����O�����<���a�@!��x�8~�Ȧ޾��*�
���* ��»��F<����{��r���>�fڀ	��Y��������#k�^����q�^��5.i}��7�M�T�����߹O	���v�_��^�)���jv⌦�lV�8W~H�_/���~�4E��qB<Ơ��`��q�SC�ji�z�p�GC����MS�Yp������yeDܵ� @�����t�9�`��+A�aZ�\8��oӽ4����љu�ՙb�t�j����%xQ"փ#�'N�(���h?0^�暎# P��A�tВ�雷.3��M��=�$���Bc��ƎUD=*������Q���o���ٔ
}&����<�t��ݻĒ�9s�KĻY�%�	�O�y_<Zy �g&&2GK�5���чڰ>|���b2LaJ&�Cd��h�s��� ��E����hc�U�j�C�ܠK��b�ۯ@3�(v��&#�̰D�ћ1���Rδ�>����G�s�ɾ�������J���])R�A���q��V������@x�T�4ڠ4��Ζ�<iG�f(�2=��龊����	A�N��� �J�ml��c�2Wg6E4;��f`Y��6�-�H��i1���KY* �cι\��� ?�	��&m�U�]3|�(-i�A�9=cTl8e��<p��}.�	�*��8Hc�<0x�G�X��ls&�����=���Iĸ�p(-n��X�)�������f@<��$�G�8��{\?�& U�L2D+��Bp�7*:�12_'�!e�Tʲ8�~S)Vְɬ�p����2�����Kn�)� ����N�ߔ �X0֩���7U��X�Z!#xb��)3���OUNiԁ���?!O(�-9����\��]������]���^b�g�ZI���o7�Re�Gl�K$��"�Fi�T`o���9�qh���8��O�{�Ӽ�_onj�1e�S�H���I�ccog���W��]�=፸����Ԓ&�Wp�� 'L���� Y�/�*��_"��I
ʠ*}�͉�8 �T{t5qnl���ſ��x������)�ˡ�������Y[U���+@e���J����s�Rghz�\w�r�\y�R��A����>ۋL��t�� 9���܆f30�:��m�R%��Y�?ZT�"?[�Ps��]F����J��
�I�{��~h)�EB���u\�^6c����	<�.�'cdT�=�	]]$�4bi�b��	��L��?�,�C`�����Oim����*�ʺei"�,��������#��������r��I��j鋺&�2qL��wH���|�j95P/��tꝤ���R��Tհ20Qi4�P���U�@Y���Ѥ�p���������*�5C�b<e�FX?8�c�Lk�rqªo����m��`ɶ{�Z� �jEӒ�(�{��\Ie��d���ٱ���7� {���;���{�����,GU�9�HĮ�X2ߖA��@t���Y�0�U��m�F����tl�A��u��TZV#��[��d;���䓿�iY�|-�����k��Js�66��-���U�
�J8�kk��6��c'�gq�)��I�BD%A�C��!�T�4���a$-<#[��r��R���#6�B�͓�^Ь�� ���|�V��-��;/��2���r��r���j_l�8���2ܘ��n"~%��
�9�{No/�~e9�)�����`P��C]����!�{�^h }��(��1]82���;*�P@'��q�S8 �,���������ӰF1C��+�sd�3K�,��\E|^ʌ�t.�O�� ��Glܫl��6Tr(7�Ou�6�*gD�I�����h�x�v����8��A8r�<�̣���s�d����Z�@�\I��k�5�<S�S9�0�Q�=^��Ð[�����(���==�ۙר�����,�4dQ���%�
e��T����^�]�UHEcJ"���C��i�p��R~�+x��<��]{޿m]u�ؿ��߿t�}?�����N)Y�>)�X~Θ�'��΁���!˒:��3�*����W9�/?�Td�0+>� ��1�A����ΣbW�Q�(h2E[��+n�-[�R��N��Ӂ�iǰ�����HM�Sʋ��Q��&b�H42VJ�d
��+N5�1�Ӂ��s�<�?�)�q
4�l`p6J�����ޓ*�:��A��F (����j�x!������n��R*r�h�,r�[o\#��2%q�
%ALY�u��AX%��"�!D�t������T1� �����;��5��؋8U�hz m����zt�m�k����X��k2�k�vh�C��:z({�ӌ���0��;c�8劁�1Q�`��y�\���؋g�X�t�H��k
�������[���'��/�N��,[t���?(��Y�tm�ȾG�3M}* ���Q|�����FZI2$�to�5�m@�|73�I�ñbC��R/�ʅ7�R=#��C�A���&�^�C��67��TT��G6�Leo �[�a�T)4X�\G�����w}���?�F�G��<g��;�{�������;+�׿_�Uk�잲 ������U]}�<���)��F5��J���63��3<~����row6<6��j�1Wf�_��>���sә2i�l"y��'f��.:���>��$G &jOtGXX�_P�UC�ŐTj-�����p��Rٰ�+�H6P��� �ӱ�C��[��W�3̤ o�ͱT`P	D�R��Ⓥ����ޭ�B0�����̙S9<7e��1y��V�|�4�mk��yy�ݩ) ���薟��
@�݁I-�u�Bx'��>��lC�I9#��AP��#`������rC&�p1t���:�|�J��*=��iIb|L<@�K��>0�4��"�4��9]�A:��@�C<��{s�3��cVY��
���Gz��5����=+닻X���^����>|�)����p��\R�)�Z?G.]]�d���X�*	'	|���˯�t� E����ʆE%��\ն��Ȍ73��!M/��O��q>�Y�w^� �!�}���x(��������JFʯ^���}�o�0�$�ǌ!�L��y�r�����������o���/>w����Ӈn^<e�w��G|�wn�\6_�̈;�����1�W�u�&P! ��ц�1S� ;)	f�=��F�r���M>Ժ��P*�+��h��Ȓ)�^�Tz-����\ P����"� �,�3\q;�  U�< 7�:���� �ce"�� j�x 㝔�0>�::��'n��G�=�l�m��Hp��eI����ɇ��W(��n��H��PeYUҖ����:ǀ�Q��Cr���,/ƁS�"�SL4�W�ʍU� <����K���P�Ac�� 1�\�ћV�cE�K�&���FK��fB�4�BK�ŀ�@p���̐�b�c��������E��[�e̠{U�����x\��xSs[P��ebu_)��M!�	�e"Ňv��3�m�M�ںJ��/�ȲRY�@��1�&ଫ���+J�b.ǬcZ�0�A�ޞz��Ĵ�Xťs=r�Vs������;Q�0ũ�  {y�]�--� �A��"��>���p��:c=������}��~��q�/���]W��������?|���=��z�-�r����_��r�T������L�H�E��%e��j����Z�;��~���H?\9�b2�+�g'�1ɘ[�#v9r�ʤ���n�^_��Ev�o��M���P��1�����>�l�׏v��rCC�#�����.rx����~���8 �_c���1��<���ER�b��i
-Y(��L���Q���d%e|��Jv�P����\N>ij<>�t���4��۳)k,�t�Q�q��F� ��M�'�2�@�=��R �4cT����+�"{�����ؿf-3���d�EXY�0M�[���U������je�����)b�X�	0%�������e_s�X�\����r!Z��@ӤP�!#�lKC��*�M�!L���+��*
Y.gl���T�F$��TL�<��5h���(	��ƅ\�a��J�ǁ������Ǟ��7����՞�����zY�����v����W9ݻ��7�~a�m[feQf��&hz�:��Hpڀ	B#��6<�i�����~�y�ER�G�vy��ν��\��J{R|	���@�CR0́YeZ��ܙ/ҍ��O�|R�6�!ܗ ���0S��'��h�Í=��E��;*'Z��ɥ��Ytk��6� ,0��Ti.V'���CM�����q?)���0�Fk�3=9�Y|c����2EY���jx!2�3��0D��u�g�ؼs���G@ů�x�4@�[�9|�D���+ӄ[����b�������i�n�&�~��=�g$�u�R$�n@��h���@�b��ew^��y�6���3�M0��@6�1��)���M��eݼ3�dO�ʇ�lHV�!�0��k���If�4�=��u���|&��twuj7����w�� �F!�Z�w���pJ�0:K��`ȧ�
x�8h�0z��)�����v�o�	���k��]������J��~�e����/_������~eƾ{%P�hZ�U�繖f�r5��{ :���6`��ps3�FS����}���L���P�BE�a�ɠ�dL �jZi�L����Ev���u	# �����oG��Җ5�-�i)��|y�e`��� <�n�b�̯5]v
M��)rH	|��g��s���ge�`?����F��^b��L-6��Y�pX	E>�Z��Q�e~m�M�ms)�������� nh�{���C�g�-�1�L,��Ȃ���8���=CLc���fM9��^����%��&�5��ߺp1��`e��H)@�[�E M�{����$�5{U���~}H��~�Z?y���?m�7��ST'FB�%�g��"6qc��z�I��+�-�7BN�N&�Oj%�}@KPu]� �ù�EX�C��̭��M���V|�����sN5,��§B���X���[R�L���/úp[��d����\���4�z�n����`<$l��$�<#��K�<_ :���)kyF��1�������"��(����>S.�٤�Ϲoo��}��	��Ҝ�(�3��YL�^����,�}�^��|�E��Q�b�Js����gS"�7�6� �a�8�r�XU��KϨ���FX��q���6��}xHx���\-'*(/�W^�'ǎ�A0�S֯]/�#s.�/����K�b䭲�ˤ�����Fp�O	HMk���	�\N7���N�v��c�(�9�u�r�L�����E��v�Z��i��l$&U�����G���8v����J�����A@O*���൒Q�&����r<��3E��5)��pY��n�h�ī�c�$oeE�=�0�G1w
���RQ$x0�N��f�m�Ҹ�Y��S �F/&�_*e�B�t�,�\uu(3�J��8�cEY�R���j��{C޹�V���D�qPj0y��--a<t��'�z�`Y:y򈔗_�/\��!��u
@�<��"�{;�XQ�����T��uw,��r.���3��]!�LA���+|�f䎡H�YrLo�љ�!�ٛ2�f!���kԊx�;�ٲo,Rǜ������-@_sӵ2�gq�f�Ub�`�޸�qMq9ؘ�>�<a���4䚁ɕ���KPtw Pn���h8h{�%E�gnj��w��~WRV&�_&ȿ%��H;Z��@��r�d���W���|[��w�r|$ %`☘.��	{�)"��R1��1h�t���t,�� ��s�É���tɼ�:u��p�;G&�+�f�:`i9ߟ.H����~;6�;�E.0�SV�t��8��i�K�a��>4-skK!�/����W�gf�&�Y���7�73��<��0+�]�\$Q�b���֬��C!'��}�[\U��~nn�Ī��xV7e�%Q.y�HB�O� ��
+}�t������)���c?B�S��QM��� ,�$����ӌ����PFހk��#����ӯ˚����w_!��{�3@%)���B����^PH��$��l��9���m7u��C�/��X�������C&�(����]rK�~�m��;�8��ZX.�\\/K�����<�R�i�,M6�t��G�ݍ����yи�3O�}���_��Y�Zj�N��.B����@��J��d�<h�%2��N�-]�y��g�`!H�પ��������G�y�)	 ����HgG7�/f���� @�J��{ &:bd��'I��H�=A=-e� Pa\�͠i��a7�p�Ï��ӭ�l/�q�V����p��`L����* ���\��[m��	���kzY��܇8&�$e��w��?z���ã3t��P���xS<ۚ+��1����!ˮ1�tp��bIGw����g�����]�+�o�Wm!1ǘn��g�D+Q{�tY�`mg��������U��/�p���au�l���k������{�{?�O}�)�[#�\]Y�T�_�VX�.g������:e��`]�7�h��('�������������Ҡ�M0dZ��6���ie*��Ď`Hw�ڒ��rkQ���h����Ηu��v�AU�S攫��Z%�͟� F-]��H^f�4T� &�����Ƣp�1-�Z�7xb�Y�sҰG7 SOO'�I�CB.��φ����^-%����~�t��Ƹs�\�c�#�����O}J	�D�2Y}�|���/�ae:�nIKMEe��9qrL�*~��%@�fٜbR8:�\y03;'w���hv��t �*I0	��hL�b�e���T����:�]�0�旤��}��ֈu`ɧquL\5N�	^m��:���s�����LD�c��aY���+&�ٖ�Z��ɥ�a�l֥0�Ա�b��S(��q��E,���2i�W��B`N98V+P�Ŕ�*���R��v �1=�k4��E�RS=�FT"J!��v��wvKgw�ڳ��o����r%,����F�*���H�9��0@�����b[������I��B����^���D�����d��׹����rኂ�@����.O�
Y�j���V,���O�-��-%8O����zA�%�ay��0�A�p]5ke��儕&���#u��R_	S=,)�
�R�(^"�z�OS��K����
^��,��CBk�݁����ҳ����Mƚ0��{D���7)?}�ϠR�z-��V�@�l�^�c]<�(�jX	�b�����t��k���E7�K)kF����2�h����5�y�ԑYHL�W��o������S"}��w��`�V�چze�L���u���h�'m��/ꁁx�b���8��"a��"�?��P�rY���Og���/Uo�F��l8cSp�Ӗ��5����
٨IԞ���~��v�;C�d�.K#)z<��\�ҕ�lҐ�?��߱A��^/��@|���2	�� ��U,�m?�h]�|�`r9Z! Ӆ�~� �Y�������g����~��;����>�_1�:=�r�����W@�l-�>����u��R�`Au���]�e���eG-��ˈ���cH�aj��m�F��
Rd�J��!E�D!Lט!�4(���
F%p�o��̰2�̛1���q|�b0�[��*�SL�l �K$��n<H�&�����~���e��n�$�ܠ�4�$Y��x�����`�:�fq
&{���C��$�o�X�O�29��3��S�w�����4�$AP6W8�B
�fGǏV�\#ø��E�hW�D;�ٴT�hm�ʲL�ڭ��y,j})2'YBňY�l<�}�d]�G�n�]�8����E�o�������lnߩ<��w����F���iJ�v����6����,ڈ"HS<Gj��Ԕ w�����˯P�]}C�J��>#���Z�pV�>��S-Aٴ�Bݻ�7(�=wVN��F����)�;.s����[ׁ	|d��\:6�6V�bsyV!�Q�;L73u۩�|+���(���*�)��-6���o�C��H.���H���z��+�W�<f�<��;��0�@�Y�1Za�ƀ�h���q�t4�h�nyx��v���X����� �0�8Rf�&��vnq�!4[/��{���Eɝ�c�21Ĥs��C��(��s"#w���b\&ۯ�tI�_Y�r������g����*y2�6gt��>� �o?zJZ�cY������a|���u����>�"�C� pL���M&���;\�8Z�y! ӈ�)ٻ��=���L
�jAC��|�r�� ����覄��uꞡ ���r�S����A;�VF-҇�����F?y�Ev�U��̮���	�M'�a�<)�{��}[��<#ȱ`�U��U��"���'>�T9d�1mR�����
epY��_�c���p���䶦V9��Ux��k~~��M.���kM� �/f��"�>�ԩ��������ԩN i��ڼUj6��X ,�+�D���0�V*h����w��)�8ԑ�V�IJm�]�&�E���b�R��ӱR9�'%?���e����{����*���N�_��Gg����\q� `�!Y��T(M7>Ƒ#�����f�d�w�ࠚ0�}�"�f���L(����F��@ݻ� T�<-K}X�U��wˬ�gH�����3�@�Ԭeyt�¥�Ю��0�X�YM3��v���J,�2���5�5j����V3k�v�fS�����*��hLo}��V���IM�7(����K�T+���g}��t������}�S��h�`〼~�O�ި��`�Et٨��,7���DsK��]4 k듲b�))�ʜJ�<l_#�>�@I�;w�}�������U���F~#�9T�H��5sT�;A��d��XMM�lܸ	n �L"w}L)�-�FN�����m ���������V�k�%�du�ᫌU!;3 i�M����!�n��j�ړ�>�A�u��3fb?�G����X� ��.��A�:σ�aOF�.�Ī���$;�/�'�x�;tM�}�^�V��G�%�̅�md�~�Ť�3n�.9��T�H�Ν��%u��`���L{Xv�D0�S��,���t\C�q��6����3��J`��;�}G2ZZ�FX�>�R�����셫'�B �)q����u`��� x:.E�F ��!\�*=V�O ҧ�TN�-f�K���Ye�=Л�Ydj�rWfƼDG�O�6�)�������յ�;�Z^%����$�~�
ʴ�и��s��@>��P��#CE<�x��'Wm��N�cf,Yb(��V��i������p�]ZJm�㲦2$[�U!��"���u���-JQ ΟƸOe5���р5�fwPiY�"�Lg�Y��c��E	)�*Օe�{�'2��t%��/J ԆZ���C��y8)ЄlI�������{?�ܕ���RdMzl�:�q��{�S*��Tװ�����5�[L��9� c��[��u��,���䀲��l�_�Ʃ��%�����"��f��sLb(EZ�T&e��]�$.��홆�)=hȯ���ڲ�Ov���6mR9lkʏLP��ݘ���^�����R
s��ʎ�)��?���~s?��Pb�.�cj#P�����9��r]e M�2���8�	2�ɠ�֓l�f͠�/KW�2N�{j�}J=��ч�p��vM��&;X�ٳ@��zX2�7���G:�2Wg��W ��|8 Á���yE5\ ��pz�Y ����ȍC�K��T&��!9��/~��`L��y�y�����Xɺ�2�֥*Zk�3�1����ج0�7e�<dǑt�8TZ�d�z5�mf �*(����U�0��*C?�h��9�)�!���g������i&n����_��{�e)[c9$#5�7��-��ԑ���BXcN� ��mt਻�E���p�˕0\@[rݷ�u&��8ɂ�oƁ������U�v��@i
��ƙ��t+����D�E]b�e޴��#�2�������|F�oϫ��+�I;����~�w�or�-m(�v'���w��2⻔���Ӻ�k���gŝ�7-`��PZM[� �\�l����Ap�!��Q����������L�Ɠ)�x� �~�R��ِt��4i0�c�6x�� ӢB��r3�@<�H⸃Ø-���6�y�}�RU� �aG��+�M�lMFY�;D��ִ��4���u��lp�X��4��
V�]�o�#��F��2�f��U���ءx�Nu����|���F�d ��������ty��p<y�;V����:���_�XP�Rk�o�C�t`��{uA�-�Ni���d��c��c���smp[� �#AΘ,j���P�~�DpsI��r�5+ ��ZP�]U!�7�*/<�\eόc
��ϘF-}�O9`��E�%�mp7:���Qnec�+7�B�;�-p� ���T'?h��/� ���d������72�l�٠"� #:�j���wъ	;��է!�Y�2�+p�j��)�պr9�_,�v���P�F�&�`�A�j�e2Cn�R-ǟ�K�xP�n��;��@ �7W����X"o�WPV�4�Z�}� ��s.Q��7�j��Vm�8'jkwʼ������E����ϔ�ʰV��&�Z���_��r��X5�^�A�8�u�8<�>s::��;	BտG���C���+��㷥��CN���t75W�/2�78<�r^\�~���[9��4,��]�/y`�q]F��A�;wإ�m���t5/���4=�:�#-O���vp<�9���6jd�l|�'%�P���1Z4���do��58OE�o3��,����5��㿙�`�|���MkژF:m�b�a1s�K�ťLe��w8�:���@x*a�!��c����I��|�y쳌�����
�r��5�gd~K�caݶn�>[����c�h�>�A��+H
�Et"jr4��NX/������c���T�Z��O�k� UV����v�ef"�2=�x��ҡ7�w��p\��?�i�Dy�UL��>��Ƞ��"���#��Q���D@Z���A�0�ezB��VY�f5�V�M�&�{�\w�����T�]%	�5����;e�Z|�{��^3�=N̕7����e�!w��k�꫶���������8���׺b���3L!�&YU�_7�&UF�G���qH"55�:>���T������籡�����F�~4��HWq��X�v����q�p�!�8#Q�4�|Rړ�%�� np����2#5�� b��ٰaYH��̜�X�4�:�;!�n�$W_�|��#r��G�0�&�Lb6s�R8ќ B�x�T��f���8�@r8$؟l��+f��T
,�`������`�a�)��QX����A�ԝ�����ͯ[y�U�����*^jX�z���i��5ç38��ٛP_N�#n�¾V9���]���9�NԒeH����r!	�2��>�f��>%��/���H�g��Gb;\���ο}7a�8L%n��qu"�# �J�VP�+���8/,I�E&C� 9�+q�cM`�9��}��Afҷ�8+��ȒJ2�uI{�\P�N.L�=Β8�h|*>33όE�a��#5dh��A*I���Y�!�@��r �Vu1jrXs����ˌ�ɇ!�޼9.�(������0�q�r��!�d;67ǳ����8�(�]��sAL���V��x��p�-����*��ŌםB��O�G�!}՜��w�l�p㭠50��������]>�s_�׋�@K�E[6�G>t7Ψ�`�ߥr���~y񇍚�3KS2RQ	�qT��B�{�=օ LZjQ�fGf����Ju�%����NY �a�Io����X�7W:�P��Y��Z�*��M�ia���}_x�GS��;�u�l���w0�Ŭ����DY�Dz����pyd�m_���ѻK�.^-_~���;E�Ck�qq��CQŧc�Q�	"؈�H�o�/�l�}ɩ��TT�ٳwJ�x�4�<�J��eN�" ��Pf�A��-@��Hw�33����!�V��Y�w+�I��=a��/��qs 8Qk"�*��&�7��F�
X�#X�$ ���e#�����T<>*הzʼ���4ͬ�		�f2+.�~M�Z.��2�����O��6 �����)E�k[0��IbI��p%���ܔ��:��b( �v���@��	��H
��ԝ��n|�X2W%��B#�N�)�� ��s6U���8,U�Z�Uޛ2�R�ٜ�rd�?�#t�^c �+��=�B!�LV���C�2���{�â��tVv����T$+�T&�M�*,��� �d�<���}L��P8$���H.�
���/źC��1L�t�����/����Z�����Z�7��té%m��>��b,�����lK�?~
��qTJ ���#����MB#x��8�CX仹�MN?�#�{h��BO���=2М��oL
�� G#�7�e�O��<��
�S�T�:�gX)(�4��r)_h3=�H���� Lyo㿞)<�M���a��HV���} W���`Sx~��I#.(i�97�q�:c�zQ�!�o깸�V(�E�3?�:QP���ȻR�֮��H���+��X�`墶��¨Y2�}�k�	4Dܒ�wb��<PЩ9u8L=.%�B=6�BC���d+�}����/��t(Pd�u�x.�Q��x�q��χ�_	6+c0F�V-�[<�5�ae�\���^��؆�gZ=]$Y�Lv���s⡥�9yh�<�JՠO�Y��a��k$S�
tUkS�E�%�sGLj�`��Yl���u=`R�L�H��5Յ.
m�����:����=�w�`0S�	���	��@eK0vO]MA�d����i[V���n�z! ���[�v�B�!]�w^��� ��ȱc��w��7�v��Bw��{��ȥrY�p���P$Pd����B]D�����J��
�h���������^�lΫI�j��X��n:#e�'Z	m�n�rd���-�,2;	tɖ���S$��(]��[��P��Yh��U�����@A�v���Vp�P�)����BY����3�����a,�����xO�1�[��J������R�/�%deE��n�op>�~qm�24�����B �O�7/Rxkj+���q��vG�����@�bv@{�/��*�.&R�� �G\�*p�� ��2�OBK���Z4��/T��U�Ǟ�:Z���2v}eU)���y�\^��FQ_W�Vq���ףo�}�b�*0�
���gֺeu�}]P���)��	�83��q`[�WImw���m��I�?�~*Kh�Bj7,I�����.%�j�wWr�xy�勤�Q��9�)�T.&
7}�k��\�:8��ܟLPh�SGNI��b�%�@K���oWʏ5T�W2�Y�jmiP��U�(t�H���pc���{9���[����e��֠?�?�0�b_1��|���`��\�ؗff�R@ԂΞ� e�}{�H���p�����G��
Y��T��e�V���_���5�zb4�==�ث� �.	�}��{=�{_�WUY>�
�z�8�E�E��s,+��4�Lw��_��Oy�a�%�ZEt�����F�����4��`�1�\_�w���z����WnǼ�"N�I��J��yo�kYۉ �1ޅd�Sn��f9�*g���6��7j��Ǫ}�l|/����z�����Z���le�B}�`�K�E� �$��� /=�(�v��Y�Pj7@,�����{/����-`����D���Ѩ`���&%�͉z] #4��i\C.X��B�oh.�tUm.��+-�fahSV����!�^��RK�=�[�td���q�
Ի��
C��?������`�Go[!`'��J	iw.���T��Uʝ��*���.[]#`En�
�O����#�.��D��ı�`e�;�0�O���N-��p� cspl������'��z��� H�N�`�gtv'湘r|���$����|���C�@l�G^9xJ܇��U�d��~be���4'y��=�vÍCm�P��X�,G��4�l����2w^�@�x�1�j���<H��wʧ� o�����s�c8�U��Pc�B�<R�Zw��l~N��oɢ�� �s@� �z�6�D�e1
�*78�2g�<b6�21l*V�|����VsY�իQ 0.�%�;���5�S�p4�Y��Ӳ@[������i��oL�Ø�A�5��	���B[����5�N0��yKB��(�ށȬ+��֭[�ۨ�e��gQ���c��{��eɗTڃإ�k����6T�|��:sZ)
Tآp�����{?�Df�E�jՉ
�x�U������᥌)�Ie����;�o�Z�֢#r(�6}Z&����a{�A��>����;�1`��g�bnF��+ �4'jih+:�][�tJ(ˇh{��&�3ƙ8!�U���?Q,��n!;�byL΄	nLp���f�l�$� F�u���ч �Πz��R7@�]�z�a1�>�~?�NJ4�����Յ�U��NՊ`*�h,I F������� �[�n3�e ����7�^�M�Xȹ��X<7U�Ko�-��e�|�:il�[j%�$ + ���! jQ��JS���g3sZ�!�G0V�?����Z����_WqF�����o��W-�fmݾMV���A(�D�jz�:,�Z��;y�f��Y �����`��O����z'I@�����/k`|��[;��������7��q>~�8�Y�?{�S^<sF����1V�a #L�0�k�a���RmY���w?J����c�Q�'3>	�|�N�%E�� Ȕ(b�̸&�%����نUX�(yD��c1�<��S��y�K���Z6��i��ˆ�R�c�l ����c���"�E(�4�"�'���(����<�{N�+]���l��|d�x�Q`U[��\��1TNef�^� �<�O_8� S k�5D�G�d2h�ʹ)aLNm̴Ԧ)$LhA��⨃v���$hyp�����g����>���]��gi�v�[�?�Fo�7��=Ay�3pS�c���.��s˵�Z;����t/i!�ʨPV����E�/@����DP~N!K��wNO�.��F��syN�9������^�:��kiy`���C�AOP�V1Е��\g�
�?/R�U�����zY<Xe��ɲl�w���_��~Ҩk����}{v���)Y����lt�*�ct ����k"s�1�T��gi��:��!c��d�j�G��O�!d��% ~r�c^�}�_�צm8� �>K\G�%�@L�@�� \���4�!��)>�,b# �@	�3>	�ׅ��ŵ	iF��_�A0̀J!�a�Q�c�ԐKp��:a�g�q�a�R1P$��kWށ��	��nqCa�u�t,<�M�bZՔ�����\��1�A�Y���W�K��8�!~�f鷒//?+-�I讼`ek�a�\���
��V����噯��)܉���py�{�h�3j�f��#���F��q�0[�,9u��젵�>� �����w�!���8�AV����q]����C�eH
�r�v��ׯ�<
����66 0�7�qctB�v�8/3��,�Ɏ�(�Mw�a#��A�	bB����tn��	C���Xa»� Q�� +��(�d
x�"��<��-t@v�z��Hhs�t �h����ka�e��%��CV�݀�1 ���ɀ_��%�����bٰ�3ܴ������ o#��{��5���p��Ԕ�^$N2ys���ι����F�Oϥ5Z���]吹x��\ǐ�6+~�<f:��c�оbp��E
E�k��j�9\C����B�$>�8��0� �/�N�`B����{�O�}�d��ܫݨ�Љ�r�)E�g�J
�AR�#�t�ƀ�qa�T5���|�,Y�@�jWȀs��	�w�?���9w��>Y���|^&vQe��ς�+	��DNZ�,N\ Xk4����E���ÃM�E�!�{�}�����-���<�@���ĥ�\�EE�K��'�6x�\.���Y�t�){\x�^��4�(�~��5�$�����A`�t� H�@�,F���`�������<$�hYb�U�e.K��YԖB� ��(�[{Gٌ��69�T�@�1�-�4�aH5$�y/�ѐ�y2ؕ���p�a��U��pG虝��O����j!9Zd��9%��$�8��� � P�����*�
���=��p�r�!�Øc�Cle�4�/����O}V�k�����?��< ����:`�sSp)d�Q*f	�]EIMk$��g!�el/\3#����|�sx���~He���V��q�e��y��s/��?˪m7���^�B;aZ�����hIc��	_�ϊ�RNܘ���#1���<�"G�F�!�|\m���W��������e�%�Y#� �d�ggn1���i?z,Rz�J�1�7���^S�`���-ǎ�y��y^��Bp� �z��;(G^> �����2Th*šQV�B�[��u��㓇�jƃD ��.����]s�����A�OaUhR;���v����!�A�z�ݹa�a#9� �ځ^��A���?0�,`y5܏��-vK4 �e���U 9�ﮀ�rÁ�A���	W��k��\>.�2Y�	�\�IX��
hbL�nI%�S>����Pg�ޜ�����=���:����0j��#XL���9�ӳ3 �p�t웶��ZC���� N7���u�Q9��<i.G:���r�F�faX>v��7��8�-�y�Q�����i�- �p�҂k6Z��^�n�oX<�v.�"�9��Ѐ��"���x8���X"�%�!�ؿHi���ExO>C�?����~o�+��Uc����@������̦�&ad�Z��lg"������K�uG�(��y�l��j��\�x>Z�I	�[V�P)��4^nzL���7#�j�[d~��P��>�Q�ۛp)"d���eh6�"�rL�)�������Q+!��P@�S.:�d�{���G�Lj����1iiO���>��:2+t̐^��*ͩw"8�-%��Vii���ܘ#��`�A��W&��8N�{���Zf����2S2�1SdNt諬;;��!�_��K�阬�<�3�&)؛���Q̯@�(��(�O��r�h�[fÙ�c��K2E��|���0o�ǔ��'O�;U��Y�&�>�ȎeZh�W`es� ���O��)#/UZ ~<(-RV��%��gV<U�
�B���$O0��ˢ�����r:p~l��;�IY8�#�믓ʊ�r���@P:{zdI�*9��]S
�7bS�4r���lH3�'��r�\�|A��3�҂x�R���F�����j��L'\K�ƣ(������54��'������o����xi}G����u��d���D��e�&"�nvz��m��&y��Wȿ��W��a���)�6��m<��� �!9͓���$kE\T��Ke�2H�U m�'<�C��2�`�VY�	�a���
�a�뒄�����M�"�RN�X��
�r]J�v^-4��Y���N9�E��f&6e���H�}V)i҄๖�v��,m0�Qte���Tc
cn-�&�Oڳ�]@��Dʾ�Nn�#��
{��/S�,,�wc�7��!d�XI�Y�Mm�lyofZi5P�8�U�SӨ�W����Ӽ�yβF~������9�*��8��^�N���ZY�j.2	Sr��Wz}1�x$� �ɬ���5D[*[�2��T�){��\Y]=&c,�+q�1U������ ��ų\J-ي��Ra�?����j ��>�A�����ʩ2���-�� #�!�&�����5(�A���(�4�|L���~[`����Nޱ���ރK���l��d=ۯ�D�y�biE�����`�BiX�R�vе5<
�0P�˙L���S�y�`��4��Z��L��;I�~ !1���˭������L�B�`��t"�Bi�̀�/��Sa�������� -\��] �Fx�L��ƅȍ�����l/���6�",(�K-�����/i���f�� �A��L���'�1��ds.�½Z
�<Z(�"C�:�_z�'eG0ދ��3�#�*B�~���=�����2�=�y3!}�{TW�����ji�ԗ��$�>��=|@x��J�¹l���Áҙ�Ss��KQ�c=c���l��f�S�U�Ǒ�
!~���|瞔���Fz������8B�u#�}f��f��$��q��c��J��#^�iǬ�|�"����p�ˊkM�p~7�p��#�Gt�"Q
>x�����[�PV�[%�.�]�| �63�T}4L�!_V�S4�.���mr�!#.�9>T"7��'�i\P�=?�.�i�z^&�"}U��/5��u��9��H#��<�Y*q���Y�6e8��-:�9��יa,>kW F�r��<�,[��`�ʸ��!�73dn���p�4v 9����L��-�@�g5w�FS��� �GL޾��T����~��V�����fA@�}M�.
Ieq�T��,�S�8,�ɮ�  ����>�tKK�t`жǚ����i��[7!k��������?b��b�U��1c�R%I�H�!�W�'S�>2�t/����#�s`¡�%���n`���]�oh�$=�H�[Mq�����۪ o����U�L�5Fw���*� |�Z���7M6�S����|0�{��T��f�K��HK�B����1k�R'(o9z�q��e���)!�3��O[u�T�H�W��)tL-�)��I��si�i*��2���I�:Dk�K��b��je��څ LyE*kk�^}<�Q���>4ʓ�!����Мc�FC�6��B<���o�a��k��+�F>�9�Ut�>�2������#x@��|�<�j����(&�Y�"c��)�u���Na 31��K�� ���-+JeӲb9��K���-a�	�yG�x�D�\z��Y�Չ�ː�Q1c���h<�=����� ��h��wv�����C��Qh��FR����K��,���U��8�}>��K�Xl.�Lm�]ڒ���a�p�	|Cp�8���hUb����K��S�0+G�=.X��2M�B]�WwT�T�G�Eu���{�f�҂���+��ԡ8���x	�A��%��Y�O����|�F�y�E�-�!�7�b�����I�$�f�AM���@u@���r(p`��2�3�n�����Ƚaʎ�3�1������X�u��,���w�%�7�L�z��(3�L�SV��*`�|ڋR2���Ȋ�����@6��b�ӟFI����R9�8�tI ����d{L/�Q�[r��f����-��s�Yb��٢�-9��>�$�k�(jz	l4]��ܤ���"�;ӊ4�q��F���U9y�_/[���h7���/y��>ј�j��U�[l(M���O�
;��~���U
���S`����L58�+b1�ۛ�;��矗�'���\=�KpU����4-Ictk%�GΏ����V)e)����c<����.�thhM����*��vU�pjY��\A(@<�R'��`�/�"+��X��>�gG�r��_�y�U
���P���R�_
	���6���|P������{��ӣd����DGX���ip`��D� `����,���$�E�7n�R�wx6�Tf�h�R�+�[�����^<�\T��'T}�r��[�a%���x�\E��E�&��18�o�T��A�YLF�5s��n_xF|]eJ;KD�R̙I,45@��ɪ���F�Z��EL����:R�B�6<3�1Dt�96وq~B<C�Z��H�15v�3�\�tu)]/�= �l5������4�Y&_��C|9�:��$�<wb��i�V����/�q/>��dנ|JGG' �q����Z���d�c�}ϥ�5�\C̎�O��2X�!�8G�������JB1@X����^��(�l�Y�Ee��]>O�Q�12�j��b��[%�o����47�O�6kt7��eK�c�Fr�qy%��ۛ��G���S��KW@vP������?�% �9>݆5�)��LP=:��Y{f��٘��ܙVQ�y�hA�b�|���Bb�V6�\*:UTz�ؠ\�5�*�/��̩��E7\-]�wJ;2��]1�5j6��\=#Wٔ�3�X��k�I��jW�<l��V�I�¤:�R9�U�W��d��K	�V{�-�)d���N.n�s5��z��.��������^���Cu����L���q�Fd�θ�!~�J����_:�}W4���Q�+�D>��`{.�)=d�W���>�)�u�t�u��a���ۍLԛ�ՉD\��ݨ�~�ͷ���%Ȭ�Y0GΨܺ��U<�(�Ŀ�a��x��s��_,K���jt��]����� N��2���XDE�U�g�{�w�r,yh�I�������32���3��|�kSAg9���}a�5��FW@���r�an�:[1'&��d�<P��Lܼc�/�>���y`Ȃ;t�i�4$Rx��f��mvZbgH!o6�~�:`i,*�v+�(΄���Pf�-1X�"i�x��I�JEG�}Cq����6�,Xk�Wμ�=ii���=����̓h�M����t~��7o��xN���)0�� ����Vq�$벖�xy�g�+YnB�D�z��d�+.%��[ˤ9Q"]��9w���s���0-y���8Q�����.�@���k��cN�mG�da��9nhr� R6���}D.+I���D,JI	H5C�k�/q�l����#��6j�v�u�UZ�J����>H3�z` LK���}yHl�a��Ư���i�{��ڥ��|��ʸ�� �O�2��/���)���"�Z9���딭�]GN&3���b&-A��q�T��T��>_�����6iH������fy��Œ
��Ed��i泲���7��\�
H`�9�)s��2?z��M��a�����(��:�Хu��VR�6c��փ�0�ܖ����d������Mf�R��=*�������2��\6��I9�y�CVG2�(�jP"4�~���d�;�Eb��}a��̯d�����b�˅�e�i&��������U��:l-�� �f�ĆW}nS������B\�bK�"	�9*$ &W#=�����R��Fm"s>��>�wf,ٶ5�S�vG׀�>������KOO�|�?%���O�����gP+Nur��S E�2����.�3�9wN�tu��g�e5#К��ok�#GOI)
b�����[|�~��R|M\���&�ޔFU?���($���YZ����{���G�6&�G]�@�5�1���̌9�����Y�3�̘��1���d,�D`�i��/�y?��'��\�r��2����kGYOW��[��?��xk[&�n�	�lQ�����\��Ѹ�s�IHʹ����`�M�_��h�̡��ڜʌ�~d��UI�����_�'�g�������}O�ܱ}��Rb�z$��m$��X(�Kj�F�X|���?�֢�k��9˰6q]��s*����G`ڀ	��h�u�Ƅ�v��B7���cw󫨜����P-AY���pI��H�ݹ6S��,��}7o���BX��gt��Q�xq�6B��z��(��<@�Ҥ3��t� �������pg�fYw�I��g�C�8�jᮃf��Mpk�g�C�V�Ԡ.5�g1������C�Bp�W~�>./�ދ̹vE�U�y�G������%��P˗o»�ʙ�^9z�� <͟W��a�Ŧ�A�I��|��Jk�$AΩbCG��H�AS���~� �3�����ǁ�a�̣	�N�;�)N"��{(&H���ی�2c������7�-&K�� ['EL:19��E� N9~u�/S�&�m6�l���������kޖM�K6�
������~S�:�(/���j�Qs��iy�`]��	50m�D���Y��diq��M�T��QZD�TY"Rj��Q)̹@&���������	h=9'�W�g�ٴ��:�x+jj�7�v�9��A)$��5��ٚ�V��8.���,e���	`��ƍ�c�"�߱̼�l<�Ⱘ8~Ӗ�"�4�c䵈%A=�H��o��8��Ų�a.��I��rٸn����#p@�"�D3SRU2���e���N��%M�����ċT����uj�����`y}��왲��~�<n�sY�3�ҳ|O�O�4�%���f�eME��!��h5��, M����N�X( 
@��\��@�6nts�F�x*k�;Ƈ{�%�ε\��i�ڎ2
��̌Y72��|���}�U��8�Α5V�O�jӢfljm��r����Q�"Y�䛼$���8æ��gnޒwVTP�DPjM�f�_���=QS��8��q2�m~E��������4X��>�������@2 ��	�̉�>�QUˊ% ��Jae�,��2���>����d�Q'�g�e6�I<7�H��H(��.�/�Ʃ�j�V��LP$�p�-AZ-�v����QF7�'� �d��I���>� H��=���=|\T���F� �x�كqi����W�4�s�|I ��^�	��O�E�s^!sV�G�����ɳ�cH1PoL�PE�Ejk��=4�^���>�kc����3]�N3��ne�t���qx��XU�� �a*�dh)3�r��ņ����JCA
�B���>�`7���9Э�s�gQ����pjF܊k���Pb��=n�)*i%��핾~d0�X1�fJ�L��\ܗg4�)�I�E����^r�̏/S��ŋn�x)%ސۦ�kW�sdS�
�X0�?P\(�;��\@��©iY�	ɢr'X�ͲY^I-�4RtQə�#���ՠ��NH̗���õ2�r�׸�\�N��W�����~$mMm������-��m#*F��m0Ȑ1�R6�j�@�Ԑ�*�� ���H����J�Cn�Al:2ٚ$|tg����}½��}�֦%�hW�Fjt����<�+s4��!@��>i	��0*�T��y�S��'��n�s7���q@�U�[��o���M��z�_�2/ԁ����K�x�v	����Ջ>��3����������vuh�0�W\,�� c�Ͱ���Y
h�vf�)P��,�� ��S���p���zf�Zy�_a�1��X�A��Z��Y���T�^R�Nb�����8@/�<s�� z<�d4�x�ey}�A���w��P@�4vc���;�رcr��?�~ �L0u��9y$���_��|���+V�0q�=��~�ߖP$�~w����ڵ+>3���j��v�7q�gR��*~�eń*	�q.����.�4��dc�D3v���^5���f`����|ֻ^���-Z��`_����d��>��Մ����qI�"�Q>!��Âio���S1�lA�%+8d1��x�e�������1t�E���ʃ?�n���'SYu�
IU�Sc-A�J�TXU�8M�G%�����;�n�@0Ɏ���E�J9��Ш��C��#�U�]���(d�&'��<Z��韧L�����v��i\0��e���py�Q�V%fpx��2 M�Ӑ���S���UKjdÒ �j��_��l܅��>�녴Զܣ,n��
J-��Yp姤���f�%���	z� )��sW��X�j]gY�c\�F0�K)/,,�� ����8��Tϴ�屗���M��ɰ�j�lM1�u}�C�����~JW�T �w�u�䏖�5b`nfF�D��K̤㸤��ǰ�9^6���m��Z[�ppU�wf��7h��UR^>G1�����W\�\�TS���`_٩��r�l;��
o��y����9ur�E[�L"p
�r��A�KA�WU�Q�{�N�U1���g�"�*�=�`5��h���q���U�C�?$3�������{��!�q�B�� �O\��b��L!w�|��b�
��_�'�*�9��qc������bY�ڃa|u��,\ᖣ{�rxO�t;	X���p˕J M�/{�;d �&�b�L5N@�H�+�����5��4(�4|��
�����5���s��.��H���K�2	��I��y�����U��A�,Vx(=�V<'�$��=�,��`Ͳ9�qm��^�P!�"���n9�|FSr�M�HYi��@�l$>#�q_ !?x�Uz�����\	ttDyB�;Ja�s�B��i+���Y#ěЂQ]:��3?Pb��H��vg�sHU�"}΋Q�x�7���?�_������I^9
~E�08Ҳ��� ��s�Wv�pO�iU�ʚ0O[�ȼ�r*�tT�D�ZH[�y�\ ���v�A]x�V52;�@����u�=�6:���mŠN��g$b��`s���F�Z��S\�Pl�O�J*�{�*����o�A��y'�=�8�
	K����B�b!V��܃Vܾ \�ݐ� Lz�q�]��,��q$G��g���F;�@ȎxԈV>2y���X���*�{
� ���(#�,�&)kU� �F�$ո��~���� ��7�3���:aj�~sh�.�Zu!������,��x���.��b1��;o�K�N���;��e`�y`�	p����B�N��,�����ڠ�>�RUJP���<���q�j�Q�X�Q�0N�v���uX:�:��`�������(������W�Tx~�|�Y^S-wܰZ#+0p�>~\����{V�v��Y2��P���u��i��d�*�B�p}�"��L,9���2L�
���c����܁��Nr9h'�Lƴ�*0���3齲\@ˈ+Q��MaR=�y7u����r���PJ�̦ ����&`��p�0��̻���������97���R�S}�ӬUM>���x�2]�f�7��t�1�(��n�ڣpo��)c���0�m���J#G:Հ��R�0�̺ri�j�J���/72�1>/����A��H�I�*2=b="`Bg3s�k5{�|���L���^�J��%g(0��V������RtƑj�{
d�l������8{��6`�,*�	�����8{��9��Wl�n8��&�g1_�~��*�,Y���2��,<�]Vl�:KP���m+R�bVY����{����X�Y{ͽ�Kc�h]1�8�XX�L�D�2CiFN�-��m�t��?����8�u�:(F<�7��^^���̆@<��U?-��Y�f���:h5�� -@QegR�z`3]��]����SA ʄ+W���6K]��d�G�u�e������d q����U<Ц\t���[Y=� +��X[C{	љ;ٟ:�1W�ۘWU��{���E!�:`�L���6�ɤ�k���`�ϡ��<Y£�³h�k�ȏ�n�0x^�;Z�y��]��]�[t:�7{�~f���50�/엃�g��5�>�8)��Q��v��eXrѱ}�[���̌��]	�,�������0h��C���Z�JM&��=�Rw�w>'���������t,Q)O @c��h��^5�&[�*U&j#�6n��j��C�F?+��Rn�܌�0� po���\��d���F��>#����@�jd0�#Xʵ�C'�vw)��mi�6�[;�h���жաh���� c����x����ֈ!f� �M�8\2�7߫p�<���{Hhw��k�F��ݞ���u�g�l	�%�<ŵ�62���e6��s�$W��vj���s���C�a0�caZܐkQ�ױ��`�Œ*FQi����^0�8 W7ݥ�l�J./l�1�#
�RT�/kb��&y�j�/5��t?�]|Wͣ9fY��0��Lr�(Hd����|KC����#�<d�Ĩ,L��kd��=�Ƽ�4=P����"�J0��3X��ծVY6,�_O�� I-���?�kn/�2�=w��{Qέ/C�`��;;��,����l�腕˖��+a�[�,1�X�-V�W��� Y3rnsP�@��G8�:�:�l�͂���b�5,)��<��
@��(|��B������x7��j��<0��*��4�����ʆ4���ӿe�w�`��P6��	�2�@���L'�a�|�~��'�uPj�������)��W�[Nv�T|3�F�YS�6����jL�	��%�%@��F �Oh���0��,���r��%UaH@��Z)�\;7�����`\�u&| �`f�+�wR�H�jT�e˖l���I��f7묷�[�-��lv�?[��4ǉ��]�,�X�PER{E�e������̛��7�E\"0�ʭ�~���p0�M���sm؊<�g��z�-��2_Y���Pv]��_a�*��T�9�RCOx`Z�����o�O��sC/�[�~"�UO���zH��͆����
{�긭@w.\�\��N��0E�ȴ�nۃ�(eh���j6�j	E�J�c�eo�5�Ĳ]����.�Z�2~���! SG�2��K�����}.ْ�ԁ��C�	����ծn̥i֢�!���y���ВAH�lI�c)��h��4(P��i7��h�B�eN�fLݖb�k���)�
�B��
ސ;��޳ߕ�O�����v�'�@�O���	��Y���|@Qc���@툹���S�B2��)�x��bl|��X��й�{p\e}��?�=����yN����<�c9��O��>�r/��ƽs�&p���k�UW�5L�F�pw��6���Ɣa���`v��%����r&��?\�'+7J6�g�;��(dMvU?7��@x:W��d�>�8N�n�w%���I({#�Y�Z�dæ�2��)A��hر��,�ʚU�!�߈�g����ıI��A�th���Q4�u�8�iu6W[��ZXs��~�^˵	NJ���熽�ٳI���ų���Nw~��YZ�b�hғ@3I"KI 0��L����#�4M���.HV�kj��/M�Z��
�� Fvj��Li��B6���o��a�M����Y��HBU�=�sS�?En>�Z;�U׹eWx1 ��h�:���YDF(�ᤚ�麡.�Mwg!`
 <i�UR�i�t���9����&�6 V��r���&C�X ��A[vߧ��Tտ������� {���HK�:�$�������rU�)?��#0+E�� K{jZ:o�; `/����a��	j���a��cȅ6�0�,�%$$���>+}����,��'�M^�0�+[�i���b���� M��
!�;Y���P���3Q��ˁB��ӿ��	��%K��"��؃]�'X��y�&�ps���Jֺد\y^�X0`�	ҏ��A)/�|`D��sǣ���R*8���P�s��A!LAI�Oް����%!�v�+C��Y� ݾc)�#wֶ�1i�=)O_<	3�W�������y�V��׊k��ucgUrR�B�d��?��������eÞ{e³W�	�<�t<<&��_���Iٷ�|��([����΄��ŀ �-Y�ɋ�A�bO�k?�s��;!�H2��=?/�m��Խ'L��1�}���yK�ޚ�����ɚ�4�0ͧ-�`�%�2��.�9u"W��R��,�g��EX�
&�p1锱�}�@:�R[��ɶ쮄�x�|�-r�C���q�_�d�CRk>Y���j�[)K��f��$��H�f�&/Z.("�΅SQ�y#��<S�EA�83�v�IBT��8vz�~9�	*�%-K���}x)���mi��Ř�o�s��h[-��?��oKgg�<}䜤^p������®ċ��i9y���^�Z6t��u�cr��!��fйۃ4(]��k��ʯ~E>�ٟ������PG-i��dX�x�� ����~imA�%7Ɣ��J۷� K#�������=<"�̴���@CHA�3J�JH<�oŲ������TNJ�U���٘�!
u.y��w����Z.�Y�I��� J���
:Ky��V��gW{
M[e�2�@�� a�aܷOּ��U^����st�_���`x��[,�!�&��:19.��68�!'R`�IB�I��)�͔f���)9�Z8��t[�WKRU	㤽 �_�a7�ƄÈ7�4!�e9�.�4�H��[�;�
�I��Mvݰ_|�	i1f|v\{u���`t�TMô5%S`��ܻ?$��?�{�c����g��lP窳0�r
ѕ�[�)Y�)���(�[Ƒz��Z��*���klppJ>��π���am��vrB��w��z�����43Zn28+c�${4&+KR3�X�2�hάp�˷=Z�d�<��\��d�1B��9NK4͓���`�Ũ�rx��^M �g�|�:�_[gN���aD$�<0�����||ˡ/�ԁZ�z�$,<Zg���Q��_�� ;ԇ�����?n޾rqH�;��u������fY�?���`BN
˺�>8fZ���q� W�l��R>?(c����Ԩ?��srb2\���k'�X�Ӟӥ^gB�2W][��R���� �$��������qV���+�Q��Iz���f����;��s�����d:4��"�I�I'e���叞I��dp<6mw�y��~N.���E����]��܏<g��£��$4� }��L�K��bu�!g�RZV�GW� /ӛ����8�B1�J+�B
��h�v~r<D���f�)umď�ݪ�h�-fj������u._b@��I߭� i���ޤ��}dƁ�<#��`_i��~\��+7<L\&�����=c?���9��h$�O<�.��/��ߏCE�E���u��(-�Nw���+\i�-0a
'&S9�h��sQ�Bh����Nv���i9s�#��t�
�b���u�BD^}fL�3P��4���q����0J7���j�v�#]غ��?�:�[���֑��׳��(���'��9�yX�C�,2���7p�d�\kEeq��	PE��X����6咽}���GC�d �-瞽 �����@�? AåA΍�;<�&��`��!w�7�����LPm+�������RSK3B��N���y����1uP�ԀnB��K��bt_l��6Uխ��D6��7#���,�u�$�5�[4+s�͟�n�kˇ�������B�ZHZpNő;nhh}���f���4IcS��A{�IʑJB�k�c���{�yX�&��������P���-5�v�{���s��tHz� �#ȻW[/�mДX� ���F�5NB�K�a�<�ͩ��2���5�Qd����s��OFG�]��8+7b�x:n��/~���&�2j0ULh���\"!p����\��SIy�p���Q:Wך)���@g�ƫ����<�(�\ǚ!G�U��H�u2~&8��+��S�\fņ�C��J[�6��qS�T�w�?{�%�p�rf����>|�y�y�nm�pʆmf���7q��A]�fBr��_7RLO�H_��֝�S��2 �b��r�O-�L��~�Tu���{�Bs-Б���l��5��$S9ǋ	7i"r"�iD��g��UE��¿:���e�	���Q΅>�G��1��9�!y�w`�~�'i��(7~���@�sI@Sn���Q��:�N�~��Iהy��Wc��֧��V~��҂������m���	���Yh_~����ߒ[�ˍ[6ɦ�u�v]=���4��.�Um  ����:y���d|lB�'\��Fa���#�ݲc~9=4�e���'er*	"�&ٳg�1���2?f���7�~�ϐ����ַzp�#�94_�>�/< �Lʫ�[����9��X�p9�]5��\)ˬ   Ͻ��,	�\�6GQ�3~�q]=�^HI�|�;��ɤ�pg�̂>�
�-H��{��#p��M�H/?=,�H )T�D(d#H3�5ׅy���#'[��i{B&��<Z�v��jr��
��u�ӏ�N޷�6�D6�'�zR���}k�Z#�<�!�uM���.�Vu��XPcJf`f�f�n"k3M� <=E���|�:�X X�(�Ν�/Y�)�o�w��_���.��m��Z��\s;Ul	^�ڹ{��u���Mhk ܨ0\<��B��̸�.�ؤ���Ɇ̢I�-0�9D�i~�h�BD�=�_宲�Q5z�9��iy�ß���n�t
����rњ�]b@M�3l����������B���� �_�F(g�w��B# ܥv/�����K}�G�%��8�l��A%����G:�`ҿ-��8�m�c�+�-��+w@��PZ�E���Y�����A���t�g���h. �501`�-�ݕ艹j̡�9|���؀��AiXw��%� ����V¤�س]n8p�?~&}�lݸY�n�pM���xU�N y�s�8,��34!(6���7�Z
��@�� �\p&%O|o����l���W��7^��/�ߦ�'�FK�
�������`]�-9t�I�&����?���747ɍ^#����_-�a�'^��p�ↆz��?,[�n�K�.H Am����wvJO�jٸa�9�/�q^F��_˘a��������88Q�t߭���;�e]G��9}Z�_���2⩮����!�T3�s)i.�`�yh����~)	��n�d�.s����Kz�7"�刺MZ%DV1F#�@S�731�ͱ�R�M׃P��n��>0�w�/�g�^������I������)�4\7k�/t��[��Ͳ:N�������Ϧ%~Np�_LRbs#�mT�����:~��rT������%��I@L�q�<w�_6�2�e�e
'��ݢ�nP����~��a>���|��P�Hp�V�ڥ�Ӈ�!�7H}cL�M���=r�|{ޕh��;����&L�(���Eۤ�>H�bJi� CfY/�U�?�U��HWO��'P|��b"^�d8E5y�k�OC��l8���<��ߐ�wWD�?���q���ɋ�65������i�J�7�T��.���(­L!c�h*�g�W�ށ��sFaSGdh�:���:eӶ63����#f�eq��ߍO�!���gkNR�i�~Jj���D�f	��F(9|��Ż����:�ၦ��%�ǩ-b7����U%�͠���Q�k����(S�̔�:m,�����.Qa�ydj�z��_ޙ�|����^���N�Jz�������3AqEʂ�ƿLM�d�� l�]��4G���Lz);͔�yl��6$Ƒ7�2u9�� ���Ddd]RUя4����v��XQr��qĕa�mr�/��γA���a�(	�p���C���[V�����à���b &�Z8x���g���H@c�>�]>oe��%���rxv�j����04g�5=A�[ߌ�Ģ��kV�ލt�[[���6,����HCp�b�~��>���'�>��`��D����[��~vf �Α�g�'���rn0�i�h��o's����1�?�c��BcJ��S�Ϩ|Jb`|2&/��|�g�+s���G��Tw=�@�Z.�w����vh��Q����'��܄c4O@�ව{�t��Q���ci���������W��� ��o�3�N��OoMR~|h~Pa�����^&!�[E��~V�;�}�<0K5y�߫�O�o�i��I4?���Ov�Km�çj���@y�~����3��ȫFO��tV�n%������ʿ�u"����G��/�[GN�Ï>��K	�sლ_��pT��F��E�ȳ�<� ���S[wl��z������U~]�AW����MWᅋ���A���`������F��`B�,V��!�{�#Ur!�(�ɀ��gfvn4s0���)�n|��� �����an�}��j���M-P?Lf�@M�h'�Ƃ�����m
1$��{��qf��{h���v���uL�3	��CM�4B���8l0��
�v�������1�	�ڎL��;�~��*�c*=����̩���o  @͌0�����l�{@^����R��v��~K9�N�z*4�F���9tF�S�˦-0#�A��V��m�'�@�V9�~�9�������]�T��p�|��y�Lp�w�V-B�%�H������`��5�"�Ž@��U2���7�앋#�c�|��b>��_K[�0b�������;�.�?'���������i��|~����4�e�R��J>��F�剩)���(/ʮH4*��C8=}�J��i�u�,g$��������[�b������5����U��R�9Rm�<0�T���R�H���gr���qP��+0�}�KW�M���r�s�s��ֳ�.�;��Q�����٢D�e&ݜ�s�:��Ks,.j�8ݖM�=�����(��X�Q�s<�o=�2/�dl���}����}�L%���/��C�I2�U�T��u�"�(`iI��@� �F�EM60�iDO�@� ���Zl��ꠒ&X��l9�J
`F��`n$�"?V-rqU-�C_�NDvlزE.�}ͺ������C���ų�i�.�N��ZK̋��R{S~��_���ǤA
�n�/���!���7�=<5��#\U��@ ���[Z�:�M�v����~8?OFL���Z�º���mh *|j�	�5�P�C�'W�FMQ��/���O�UBP�h�4�K���d8�8uVz���o�]�5�3h�-�I���Q8���#��D��G�Nn�����~���Yd�ٴi��5����HD~����Fx�z�~ikm���\mrv^M�����)�iz������Pی~(�?�j+��g�M��a�Y��?��<)M��U��(\f�ʁH�nX߫�X�+)w�����['�Ĕ�xf$ `���ۯzb�MIL�	��y����R��L���t�u�Kb�0��̕K�(�Ƈ6��V\��)ú��s���'Yj� ���%��8���w�`IE>�'X��)ƾ� ��:�5�e�,O���D
��v8��حy���� I����G������=�̓�+R���=QHV���;v��*&ɑ�%�v�,��?DC~NM1B�!DC+�2��,"?7��B�ᴲ	3�����Q,w�i\�P�ER.�GM�dB�4��_�F/^ �[@���Ur��wZZ$s��S+o�����8(��zD"�9|;�"*�;9'�qL>��:�������N�NA�4<�򽨏�����f09�(a�	&*t�9�VcXn��z=D+��al��"���2��`��*���"o�B(>�瘣+>u���e<b1 �<W5Q6p��RO�p5p`�R�f;u�U�v�ښ���Y~M`Qu���9nx�+˖�t��B��3���n�S�L/�hs�9���������dln6�I�z7���A��c���R�g@O�5 '�L3�
�K��ėxn-���^��B�*�������Ҋl��ܼvT�M��/��'i*,�/�����RM���c�&��c'����3�gߍ�����d��w@�ƠJ���?�/�]��P�C"��y��ɚQ8�S��U��+Y��� ��ˢU3r�#���9|y�
�� �y�VB�_m4�����h��}$����{OI����G6o�_H�Is�1�6���&��"���%ǜ�!2*	CE�-7��ޯ~�CC �IiA����㕭iB�6��3�4�RV�M��b\e1�!��C:��}~i�v���<+!�4�5Ț�K�?(R9\]s5_�:*jX�Tt�j!L.D��t�i����a	��# � r�^�*x"���I�<R�`�#�	�q�]�~Wݜ��V���v��Z�k)RY^o�ss0��K$?��i�����& J�Y���ŀ�5�a�K�=s�Z�� kA|8'oJ������+�F;=W��$:11#c�f���Q����%�m�KwnT����Kh��Q�oɇ�N��q��Z5���X ^@�������
h����+�_-u��Bӡ��z'u<��_55m�3`�v~ͽ�T$M�4��4��E4�b����^D�N�'(\�v.���9��·��q�,���|uKu���ӘS`��W�O��
~b9�����sF)U�N�-��e]ؿ�'go����y,4����J�u=�G(7�e0[n-\���X�ϒ&NkÏ��f��9P��!� �ٖ�R	218�z�qprd< �8��W��^h���v�n������/�g���8V�8�)X�30v"���5�:#A�anH�8��Oi��x1`<�xTU�R�&�<W��A�Jϖē��k�kg1uD�0�����kt�6�Qc���Tm����eI�K?�p���,��G���u�����4hJ�ʃP���%*&8�	��12�����::�Y1�ʡ�ʭ:�N��I	�_���Kԭ�k��S�����ȥ���L��q�s!�b�X�1�]��UYӫD5y����c�'8�!/�@U� �e໴|�x�j�b����\W�l�ń?&��/5Y��LT%ϟp�0��a-#�������u�BjHj��f�0CF���u�u�"��z5��&5;`��:�~J*�K	�El�ʣL��9��L��i�8���t�&]~�ը7��ٰ<uxH���a�0Q4�5F9����n��r�	�!c������@�"5��-���3��<�$ ��s޲��Z;�K��n�=�~�0-,Uau,Q����Kn�W<��_��C�3�7�geݙ#�N��B}�cbYph���E��	���\xȈ�*@ƹ �@��@�>���v\�+����f�x^�`���Řue�����F`���-� Z�T�-��]�..�q�lpb����i�M_���7
�|��>Il�ܣ?����W�,S^���Wsl�	�1�-��&�5�$���X⼌N���W'%��TC�c���l�U�W����1�U�yZj�x�U^,.�|�o��_uN�N���$7��˃��p�Q����.t�}��!�%f�\�AX�A��Tφ[�q�
��hPjm	@�1s�c�0�]Zu�.>��j��A���ʑ�2���W�[5k�͈n��bCUm�%�.s�}�1E��2���1�S����F���w�����mj�W	�_��ST�Z}�psu){���<���j�r���7�r�ɲ%�<�p�*q��s��P@��GJ�
�7~�sFz3044�,�n+O��t�b��UJ����G�tp�x�I��<��gu��)��另�G
(�%>��=a#<���"�w����t�i�I�a��4U�Cx9�)�w���aRQ8��gS�4��������pL�fp��as8h������	��]�ŃFm�cQo���G��{.;��Wr�e�d�Еv�����p>x�^ٶu���h�F�k��cݥ�Qy��8�t���:�)0�ιԘ�5�K���[�f`_x��	l�rvy����dtn0�j
Mi�3���%���I��wK��H��U&�9#�;�r���Q�O0=Ƥ�l,S�X�*cKUj!�g�=3�"�����7㳤N��$物QP%�$a-����f�B-���S���5�Ww�^��{�a�3rա#�Q�4#�H�h1�)~��a:�b˟&� �{�4xs1FHb�}j�3�C#O�|�����̥8�yVI�,�*~�g1��Y���Ԅ���M��u��w���&`�a���iIE��-(�B��,��v�Y IBX�^�)Xvlv�Ɔ:���}r�m�L���Xő��յr�b/\D2t�,�	"���\�H��I��"`n�%23(��S��:D47�*��Vam�M)�(�f/�Ϟ����n��k�=[lp/@E��Mu9/wMe��ʞ��o�R�]0`B�+�ċ�i�������i�f�W
�<��\̦�Ck��mL_gm���.Б��)��@�PP�OF�6�5
T�!>�?�D�Y��#2�ۛd���$���nl��76���T������>��ɍ�`��+�g�}vj;�,ͪ���>a�	�i5��T���z��]��p^�Pr|`���I��Q�#�vT�u����ɗ�F�!����B x�k�*}��s��\�����r��$@�9�A�Zh%����Qy��QjV����>��ޜ��T����,�6�`���S������ٖf���=��V��y-�s���;e������L����T(��}�r���j����km��r��?�	D�=v�[�]�����jG�秋b��n��7��G�о$k?31"9^֝PF匄����&�@����q|�љ�Ƕ�Sh��?�&4�FLG�(ʧ�D� ��P* ��W���}����R�S�d��g���T��f�.�Q�DM��w�{n�Q�0q���Q�T�շm�������4򪽖����>�F-�C�CB;��Pd��d�3�_ÿ�}��m���� ���[b�I4]�w�G���r��A��m��e�6����*4����1 �0W�n��`���=�
�47�5�CX;��193��ӌ��Ȁ M����Ű�̧��g���33R�#}i��:�+*�C0��	�Uwn������n�Ï8
� �M���MN���y���v���hW4���ɪ��j��ZO?�a9i�A:)� k�H�I�4�0=х�:ټm��=�8duR�{�e$��BiT2�ad&�.�?��a%7/0a�ȉ!���� ��u�8�s�jbS���MF��"鮗	��9�b����}0�FZ@G�ĀP1ӗ�B��3����ا6�ʩ���.z�sh�t�E[�3ډ��i�:,h�l4�ڬ.�'��*P�!YU�i!7[�M��J{���
�Я0;���&k��Lו�,=�m��ֵ��@�-��n������|c�ۜ���S�ZC
�8�R�K:"�{�K�?�5H��}��rt�$�񁾡��+2�[/�V(a��Lxos�G�Z�ʼmε� ́�3������u43_�A�!�����Kw�>��Ƭd�9}�~i��*�����˺�3���)�~7s&�&��^w�VW�^�����Bz���R�R
z����F�L�Vy~�ܢ��5��pŜ�g�CөMe:�0���^��)��=W���&4;.�AvC���r7�E��2|28+7����jj�o��_������C+E���;�;�Ŷ]n�i�L���n�4���Xs��!� �ǃ�8�(���+5��N�]0`ʳg\���,S��LFS#���"�UQi��潵6C��UH��bL�>���$>�ŧZ0��� 3
�@<j�l|H,�Ir�Ylx��,�y���z�� ��!�l�ƭ��Ƅ���Hn�<	��p��h�Vp�$���l����&�/�7�$����Dj��]
م���c"��фWj�Щ�b�8���ҢZ2Z��n�/T��K�U+�0���
C�� �DUY���ŏ0���_�Q0�څ}BF�2u���U-��1�令���8j)��䣪e�`�T���������CP�L&"�Y�Cy�՜�9�[�	Е�����[�y}��bi�����@�r�����/��$AN������o���>,��;����e�S�Ÿ��s���I] �o����)8����hi����k��
�f�:qN	��S���
�{��sZ�������dr)8��e��C�ʶ�ӺEl���8��`޺v����,o=���#r�m�K]�:��<̣H�:I$��ѸK�>��گ5�mJ�\�|���L�����G����U���ݟ�i�M
�]��Ř4��3��D��d'q�"��s�?&���4��wuO��a�s�y�q�;��n;������C/�ʙ�5+q�������h@Ά�<` Js A
7P�'���h�!w�ϒ:xW(��Đ̘�Pv��bj���*߭�1i �j_\�8� W�'�|v���j䆻��B:��~�<[HA��6!�DBe�8�@�c)���[��L3��U����o�d�����RKH �~Y<�Y�r�PX�3҈�����2�ڹ���iSS���`Q�j��'i�>�-��D�>uv���m	c5�x��Uؠ ��i\t�1�e.Կ��g��k��d4�u�o��L�Ⱥ��sƇ��Ŷ��M�1��w�p[-F��G��Hd2�}Df�&����/�=u�٭�����a��!e��
^�eB?�P0��6aiki@�k9��hj���6	�svg�'A@�	�-��tG:P��K?�483��~$ׄ��wZ��1�)S5"2�;Ǟ�Ԉ���j5 ��j�-%��%_������qy×�U�?)ֽ[dݭ2:ͺv���"A�-!�QHւ3��h4"DFϟP���Y����ى��qoy�+8��W_�����y��@�c���;0";׶�7��z9   IDATV�֯��M�i�. @��LR"�Q�D�m�Nٰ����R"Ȫ��G�˦K�2�d�� �M�p���	V�/���4������*)��" #U7��P �Bj�=�ٽ�fE��i�m�6)�_�#�K�H8s��oLɝ�d�|�����ᢍ�D����m$"��b^���@c���lM��xIl`bo�*�i��5�c|w�Χ	�Y�'̩gb�qRvnΦ�6Qk���ݟz�54�;�3�.�aڧ[�3$���(���q�R-�[�,Z�{�'k�rww�|��a<�;�Lj�>x�QN�W㵓C�P��^�s��)��܆D�;փ�������2P���err̘�:[�5/S�Ьb�6�X�D�k��vy�񧡝�$�-]�+{�F3���4�^�5�;���>��L���[`�3��Y8��yߝ������Ԧ(Z�"̱�=Nc�8@Y��Z	�����I��*�y�e>&���)M������܈ %�	�����R����hR���)�;�>S�jd��<k9 -m�T����V�I�9�&��W��6yb��e~5 ���K>�܆�\��t+�l�v<	�J��0[�mnȱ,�ΐ����GS-�S��yNv�]#]�c�FZ�\aȓ�3*���Z��:ӂ���H������s�R����_�'�)���s
Ѭ�+D��Q���/D5�9���z-r�_B�Eh��9��94Q3�յ��T%��n��UƉ�`�w{�� �|�@��JG���M�4��64�ISG�x^8.��#ҍ��P�Q�p�Тv%qXb��OY�3�M�=9]�UEchv��2N�N���:�1&�9�y�i�͠|l:�Ϫ���_%���@:���;���h4����52c��6&\R��gW�5z4�pna�P׊K��QKWk�e�5f�D�}����%�0���Ԁ����[�������/a�{e󺵲q��Y��F �2����Gm��#������U7���!_8p�`�&��3��bXk�#���ľ�g���>�������3�&�S��>ML����a��=d���M�m��?N�Gzz0"o�a����B�j0�e�w��t����XC� �B���~��yi��7�����[�xd
�x�ضs�$�l=L��R�몛�˳�L��tg*�I�L:Ny͉��tQ�v)�v���ĉA��n� K�K�?"������A}m�V��{�W�%��Z��٧��u3ҟ��D5!��s�7)S2o���f��7KS.�fA��9rJ�Z�fy=��Q���'0�'�`��	J}�Z��̂mҼgҒ�ה�s���Hgg47qP�837�*~�[o��~L��g��樼<0&UF�T ��Sh	p��V�&��Sq8�������';���nA˨�'�S@ftԥ��/���[�q4��g��.����g/�����⩉x���L�DJJ
�vl���#�C��X�c8A��]h� ������s8Yf�[�+"�q��u� ��9j^��G�_W'k�t�<M;@Yp��`���[I�;�R�D#�G�#/e#@�_�E�5?4���װ���F�՗�_�+r㾝�@ta.�@�@� DJM��<�Ղż����!�-t�}}9n�:�A����'O�&�޾G@`�;��;x蔼y��M��4�YW���N��}d<U4�C�ĚLMJ�/�3�L�C����{/�V����D7�k�4S�ތ5 �ż���i�#�6eM�˵�8���v˖��zȵm��K��%ە|r�m��k����O��>}�p8���?��əG���(Bs�O��_�M�X$]����ڱ���	utB�2�\FMR�S( M������'�%x�H�<ur>�_Z�c��c�G�p��0r���<[��td5UM�>�N�پ5vk���J��ӕ�SY8��Ƽ�b$m�9T��<���Y���ӓ�3����̌������Qy�=�Ɖ�!��U�}'�]s{���:�﫧�\� ��8�a)$눣��*٣��� �j�5i'����L�$��kg \�)��!��[w6����� NL6oj����������-lz&Y����̫It҉��r��7ʧ�W��T/o>%�/���y�N}j��]Jɏ_��
3ϡˉ�y�e���zc#Y�ǖ�4�QS��v����fK���AW�ó�ʣSy��Kы��#˲l�3���Ac �5z��)�x�Ac"�������W�o��}|�B�T>��ɳ}�hؔށ1��Q�
	P|�ݒ�|��Q�K�����}�hR��,�e�ϫ�3�5|f�^�Ly��'�?���a���Yh��9�8�&`��������h4�˱�Z)h�/�tȪ���vF /������v�S���[��V��?�����o�L�R��	��:������EI뚜�؎�x�	/�ZYV(�NT<�'::�|*Xf�[�G��C���"sBF�h�ve׊��;}ڂ�Y{ޫ{zn'e�t饝@F��3�d�׺�ޮ����Ʌ��I��{{��ѣ���}W��'�����x���}LiSk3~�$>'�����+��ӷ�6�1��>@ͫ�0k�J�Ʃ�߶:)�Z��G�Z^X's�? L�p��D��+�q<9��A���[�t�l�+5R5]q���}$]4�c�0����Qj��Q�fҘ�����T7�������S~�Vs��(�x�Z�E��[�P�'��U.���m���3c<�*j��֐K�PQ'��IƉ�J*���v�g����6Tr	���pZ��I=�R���,��bG�s�m�^<p�D�6�.�J� ��o�k�y>����.���2�����HJ��c�!T��+���K~e���AW)j��'�[�b/�L����������YN�n���`��K�B�pĳo��!f��^���Y�3l^�}�|��M���i����C$̄v	�JQн���r��W@Z~��^~�׾l"�r�O@���}�����5e�4�M7��u�Ï� F�y�f����<���{O<�`����O˶�Ʌ�&���̎n�ه�����J݃��8�1�=�d�15�II>���e*0ȯ��8�&������LU!��*v�o�$ˈEG��+���q�5,�ΒJŠ� e�"; QE��dk�Y��D|�plVxi�'f�`�BD��N�ns�!����bltR�8D7!�22P�����X[߶Y}�ܷ�Ԭ]��u�S���a���;b,�˯�#Э\�� ��6Nf�oQu�֢scf� �u�jZʁ��0,�}�/�g_Ӄ��]/ȇ~�����6�����,-����+?*�X��x#��Z��+�#�^x��������765��ג�n��N�nzm1@�rx�b��<�����w4~F��Y��ٳ
����|AG��Ab���{$���������1��B��,��	��8���#2���;emCTz���7�"z<�?�Y(�x7
��0��MQ�J.� �G���Q*��0I�q���hq��R��A4�X�_�
(tr��։��?����Ok�|\�`���w���}m����K�_/g
���v�2u|x�u�k�!����Q;�p�L�~h����\������ �@k�Jd��£�������4�im1�����;���a� �6I��I�6���������m��5�lJ��sq�|3W!�ϑ>X����n���w Ŀ�>Y�r���jڪ���Z}��A����F [DM���4�n�o^�c!=�L��rpg]]`��� �=Ԟ�ݠRq�ޅ�!��i���,���eTq�,�����a �|����P\-O�붮YJ��5s�ߣ_@��d��9��o�#Aα�%�MKKK����[r�����<�'���Y�X2W�o)4��(:\��*�E���D���|>����s��0��aT.=�;�ԛ�a��������/!��`�D�M���ظ<��s�R�0*�\8���{���!�[�(�=}�����3��_�p͍�r�[�XP�f������3|
Ē�3ܲ��X}}Z���0<��qm�m����,�q��� "�o�h��|_��m��4�q���e���8��Dj��ٶ �ql�j�#?��G^8{�}���~o�d��oW�]��φF���?�rj�FX�=11!�CC`���;�6H���C���2��4���T�p��m�(�W�,�.ǎWrcR
hV�`Rb�E؇47��4}vԃ7اN�N�6(u����.�����@F�t���}~�Ċ��� ���m=ɚz��&�=g1fi�3*�O^ X��*���Ej�b'�ҧv�`� <y�2e;V;�m������ ��E&k�ɬo�lh�ȝwމ��<��BhM��!�<���4,�npl[*���R#��&~k|W�g���I�۔ڼ���2p��;�_���Gvl�)Ǉ���7@] L�FN�"�g����ӣmc[G����YN	K-Qss�l���ٮ��5::�3��~�	�����Y��~Y��}���A��N�I�zJǽ1bse��芮��(�hf�!�D*��#D����s���[o������C�����+�-&���z	��ߩS��_����(OS�=j[|`Ϯd-V��+tgYZ���|U���~Qn��&��<P(�0�������#j&���}�u���!k��@��ֶ5���i_�?^<��[�M�����x�G���>�F֭]#G��m�^Z���| ��l^�e��Lw�);�yr�����M�{��ߗ�5I������;Ez�;V@���.^�3D5LG���Ͽ�_��$/�E��]p���(��x�Z�\������w��
۲�>0 ��>�gn"�S<�
��jp�����
�)���hZ���.���t�����ysVƦ=2^�"�~�JK�<����jF�B��PU��,|�,�B<�:�&w�S'���;�e���a>����I�{�~�f����+�Ι�����Q�s��i�Yy��;�=~Z>�O�	�o�¸��X1β�����]�m�*�Ff�^�));@ഩ���{gg��Yg6v�ޔ�oZ\�BXꆲڴׯY�ZZ[:�lg4����{���g�]y�0E(���.0�+�-G}[�bW��c�j%��zC�+�Q4{(C�sPt��Y��m��^��E���_�w�|��_��~<��!ujnkCԨ (�,t!}ef=O ��͓�=a=��S�*b��4AV�+��Y_�!�G��u �����M;�,�+�k?_�8�P;�&uI٥
���{�����Jca_�>&�:�����_/@�4�ލ��G#��~�t��A�������:��T!+ �UYt���ĥ�kٓ���y��<���������Z��6΂~gwې|����̹A��}�Ȁ��{n����������[��;gZ/��𶯂�0�:sz��v֒X����:O?V��[�Z4���U
<u�d�T�H��A�+����0*���<ʶ�kkk�	��#�*'ţ�:�Z�U0��F�}�]F���Lq�y�����6�P�9�TN�8��G�{�{[SQ���y��Y�q�sIW0��ɩ �pf�$�"~If�}�G�B-%S�7�155t��ϳ�Q��ֽE6TeU��P�xr�)��X��
����`"M��4G� e�������)/��T�#ذQ��VD(b<��N�[-('�A�P��i��:ƶ�ZcN �6:h[f�>M�Qx~e"ޔ��6g��@"t�A�QU��T����i����Z�<a���#s����6YU�q��`Ԩ�m<p���wA�;�N"$=m����I����B��� �o���z	6&CH=4E?d� �V��A���)@!D��J�a�s�(RK�0�4�B<�8�t�!�!SN�{�R6��t2�i�M��&�FW�`6@�L�[P>?����g���������Ø	��_��w�Sy�Y����1㐱w�v����V�p��������_��v;�L����;��f_��|�_X�
���l��O���H&�*7�KŪ^���%�D�Y��z\�{���g}��}�6���̧I���~
%j��o�&�����L�O��d��)y��y|�@����F��T����7�Ē�P��(hҍ��u L���hl�JwdU��C��2R;t{s��??$G��ʸt�u�G>� 6t4<sr�B�B#p��w�����>��l��'/@�zdbl�9]F��Ϋ�����^������4M�����Krf�1�E��j���|�1	�_���U���U�`Yڇ~����" T�Z���5�$:�1�G�b�=�'�铡��7C�ibL��~��_ӭ��6�Ћ/��o��i��ݏ6�D��(�:�����1&�D���$��)ȴ����4F|'7�qp��Y,�K%Y�il^�x�Z�<��T���c|�]��Wc����ї��ofc�*Zm�<���cdf�z�����~$�4,Kվ��\>�@����rp�#O���f=9�ۚ`�gH{2h�N��õ:/5��?�m�s��-���v�#=hT�'�J�Fr+��NS^Е��	W6�<݅zΗ�����w�]�"a��oE>�R���\{��M?�C!"d�6J��$:�@&_M�&��R�45=�	l��vD���$�y�*�kE3��=��eO${#������7�i!]�߃�e)f0+�"�5��N�����1 �@������_B.����Z�0���4�5��R�V^2@�����/��@��aF��,��i�
3��F�Bh��`�����������p�����7�)鯂�2��q��l�t�%�Eg��xs�	��H�`MB�qb���/B�c���x�X�	ʊ�*f�A��&�?�:>zLۢ�VEn��co~O&��>�Jur�9�/�$����0d�Z����
~��
��'�I�.3�"����cC����tfd��Ͼ��%h������$i��}��+6R
�w~B+�n2&T1�sN���r������fˇyx����Q�`٢��ж��̭�iϳV��~A�����㆙i�3a�<Wm��4���g�׸�"s)�h_�="_��yQya���uՖ;�y�g�����s��ck�c��?���� LqԮ��ζQ�C>Ϥ�K)N}j��9+'enO�4��������܃`�����%t�N�'��_�[�q0�i��Ɨ)�PK���A�ڵG����J�9�y���������b��ϓ���kr��B{l����I&;>-�S��J���B:��<���&0;o�ö�v~,բ4q��ts̺��fcWb��.F����݉�\V�\�R>0�trv�T��Qʺ8�s�$��<�YP�z�x�"H�FaZ��n�����сQ9Bh:#�	8�����
5����AgX�i��9�jf�S���g�'J��F���H��>|>�U9�[I��Ҩ�qi8$���Sz/��z
4|2	OO�T,���J+��� ��Ee��+=����?3�G�w�?��a^y1�L�ڤL^:$�?�Ă����5��8��3�d@e��M�����:�k?ӑ�/���wٲ��x�r�q�X�	�H�ֻ(�*^�K/ �f�:�<���BP�Q�.%7th��az������l�9�}{m�6g6���t �\�����>@ )6M�댠�z�W{�����~�װ��<����)J��v�����*�����A�>�>h3��l �K��ʱ��_y=��x�d7b�L���>��A�@OSv�x�Z�?���-�n�����w>$-]�EJ���W��
�n�Dj�l}�_����t��y���q�jk;1����`셟=/���~T�Z��Z�rǢ��K�ɕ>w�݇L�(P+o��",6�[�<�k%*��c+i��]ޓ���/Sf�{hYW]�PcP�/�U�b��Wfjr
e:W}< h#p�>��q���92]�b�Q��)|A�?�nM�:�L����oJ�y�$�,���sPU׺�t
6�0m"�7).��d6��H3�7�:Ʒ������j����b7@��W7�Z�5�Z܈���r��Ծ��çc��`U��E����&F(e6�Jޜ�n��R�n��J^�\�4SXZG�^-�T�O��ѐ.U��F��~���&�E͐O.�nͫ�Jc��1�Q�Σ�Q�T_��@Zx&��]��@a�pA��6�u���|���a���:R�G@�38�ٞ�I�$��k��&����i7�k>�-�/^5��y�)�Z����G\���^'�C8e�mvS��u�R�EIrjq��QbJ��1����o@��wH*��D���ɫ�C�ҬO���r냟����28�Ca���HlN��p¼� }S1��v�#v�}�ș��F`���DٗM⻐~]��h���.�/�}Z*�|ौg���u���2z��K0�TyvK����9����6�qh���#3��]�,Q����
��Ū25ܠizcĜ�(�l"�_8ڎ�6���@`ǦX���I���0��'vK��l��b�R��+����3���T��J�1�7��v5��1TR? �u�qy��Q0��@I��&d�h���i]5MˡX�Z#��@-G_��>c�j~I�G�J�<>����{�F�8�M#���ǂN-��:t�!���jj*1�FꐳPM��.Q��u���}l���+R�#�	;w]����*j������r�BM��7�C�k�k��Ҭ��i�������B�w��:��`���,�	��L�������i��Q���Íj���U8h]�a���*Cć'r�=���_�- $&+v��*��	Y#��[H��&.���čVO�* �H< �=k��Z��j	lz�����4O�JY��UlW��h,�IJW���d��2�s���W΅<��w!�W�"���\�t��n�fC�����'��2*�����Y+L�}k�L�Q�IU��TPc���MO��ɱO����l@�	�ZnV��n{��0w#ެ+$t:,P��� �8���*�Pt&�!M�f:_�a�k@�s�ݸܲ�_����	��a�xD�?��Mp	kCtܔT��QP4kѯ	@}i�[����I>�Tl�Fn~t�����;���6.�ܾW��{�|��ߗ7='�g^����ځu��͘s���c��yѨE<�`���y$��7Nm(D���o�(0lR ��iP��[�=ۥĆ�&8�X�������Ϭ>�F,I-��h��ZMR�T�ހ�cSO�l^�,O�ޫ��>jz8���9t` z�Ue�=N��z�XQ���gJ�e����(�~g��M�q>���p��=�����!5�mC�6�p��<���/I[�'��&��
XZ��s{;���
��~$q����n�r��ࢮ�pA��fo��Q��C/��M�	 \�I���8�U�f�Q��ः'��.��k�_����ޖps�­B}2*��Ԃ�沣��z�F@�h`M��Ut�6����+��ԣ�#k��Ț�keI������x�O��_�>���C�%�{P����o������n�[=r������20{���x`*��� ����6,乤�Y�&?��wK#o��Ny��'��|X�z���؛���h)�B�����F�3Kx�Ҁ�)8��o�ў�f�sh�|��c9��(�O�7 |7�y���^����{���}�MͲ��N�|m ~3K�!���S0L�4U�k��p�O㠷��nL�KF�TN��[�i���/����+_���8L����)+�P+�5�T�2I{%�N�(v�F
��kY�]���L5O8��y~�ӟ��{��@��K+=��z���j �|Fkg)�.My������J�Óh�p��!d��!牜�#ɰ_мas-�^c}( ����Wy�r�"_��jZFO|W6l�%��_~G���D���{�ȫ��U�[���za�i���ftI>�K�Tn��@��{�]/s?yY��y��X�_�P�2� �iF���[V����/�h���ٚ��6&��$�Mߎu=�n]�4<x�<."�0�V�HRDLd0�OKO�$u�1\H��q�V���q�����V�ӄ�jV�O�l.��ͥ:!]�U�%
�`^e�O���]$l�I��~J��%w�Bq�;o�V�����7ɻn^-��;/��$��)�Pk8L�]�z�<�v��JDi�%=àߨ��!hC{�GFqѿ�����U�-� ����_ڣ5�����˞��#3u7�\�0�d�#��N���vV��˵s����B�����Y,�+�P\�]�v�z.w�|�EmI��&�\"D|�l�)������t�@Sm0+����>5�]˅�x����"���#E
˙��^����L��Y��9p����}]���AA]S߁9�4f*���s��\�D�-9�?�8?��s�1�	�D_7n�����gec�L9�\�	�MC����<���a��f��ݟ�O<�^�������7�)�?�%�{?!�c5Mj4���ʳ�w��QkI�3�����B1��|0�Q��,$`M��\�t&�F��]���i@��0�,2T�G����i��4g*[��V0m	5a��hd�Xc���`\�p}�1��i2�	��Ir��U	 H��G$������e�g{�ra�Mn����;�5յ]�#Ȅ�H�hNy�Z1u�w�#+�]��3���{ ��58Zo�6/`��{�@��G���l�ckX�=�6���8������,u���NVuf� �#M?�%^��m)���VK��Fh!�F%Sbب�%�9j��C+�ߞR�4Y����F�羯�Ɓ>i�G}�΍�t	g��օALk�jÙ��UeB�	���J����׷Ȧm��#��+���/�����нȪ����phՊ��֌mj@x�H�sy٤��^�T-0��Y�����Wv8�Ԃ���m=8��̝����ypm�xh��/7�[5�A��w<3�f��x�^�9"�l��������D��*���ce9�a����?*g�D���M7����� �Le��r�P�y:$Z�3�3��ju�^x�;�f?����,4�����Wo�	�{@��'���]�^������p)���X�M��Y��>=e�����T��!H������nt��Vm��Q����'Nxeb��Ny��`iN������Na�SO'd��Fim�F��6N\���H7c��3�7{��Hl�.E�+^�E�{�����@K�Q�p�� >
3��|[J�������Z��	 d;�k�yތ�Z&j�HMn�Y&��9y�y���[�~�|�}9}���|��`�N�iͽL�Lz�.8�C�B���K�� Z5��R8ͦ�2���$6�/�n�OR[A:"� zE���!�/LJ���x6�ݩ���~[�� &y�m=����Ӂ�S%�%��h���r��3�`��j4�`�sz'�"�����B���K��6�����yM;2kx�I����x1�����A���w�.i��n�d���y�b�u��W�����ƙj!ǀ��]P\�ה�j=_CT�c~l鮑wnE
	���b©Ζ�.�O}]����)��E-�L漞�[S�v������'��¹��va��Gsl0��TI-�H�~O��\�)lJ���1�`�vjn�	l�
T�]�s����m����t1*��� ������y ���=�3��H��33Y�� 00��>=��ID�A����!�ɟ��N�6H�u�� �H��V��v�wq�	ʊ>C@����@���$���_)N�,8�k��d2'8�-<41Z���m����XD���ߔ����������^#�5|�p�!�d�@������j�׎��d��ېیO�F���1��T	U0����f�$�������Q��n����ZY2���y�}r������c5�"_�i���v1*|�����[���Bc��sJ���ߗ3�.j}ǎ�X���_|��G�y���-���.��}+���/��"��l1�[��V4��ݣy�g� =���������G�R����g`bB�G���uB"ѳ�8������8|fQ�BΘZ{�4�rC�\v���͖�����j/��ap;jI~A}�|���Ih
��ġ���"5m�γ(Q$�� K���W�>hs<v�?�M�#�����W�Fn2�@ML�y�,T-AH�rj r����d�w��ѝ�l���j0Ƀ�"�"�y$�d*��`���O��6���ј���Cs��Z;�`
$���=y�X��jZ`blks.4y�k��K�x�	 �DҟP ����>�`���J��ޱA�?�_Lb���|��.=�l�Ɔ��sJ��Y2&/r�5���v�6<��<�7?B��z�u�ߕHÝ�	��)?�/d6Qi�,0��K ��ƭ z���<�d��*���#��� ��Gv�X/���q����9.I�
u���`����ؓ�'����F�)�nۿW��y�?��07z��$�N�$�cb����y�5������ܽ���Т}���>L<�VLr�ֱWՃ��7�8�nc�@qS��%wܩ�v�y�j�9�-"M(��u7�ʚ�i�N�����%�j7J�ɸ��i����2��s��ѐ	ܑ�� ��w~���G~��-��TE��!Mo�S�"`��U�����!*(Y�|{ؘ�g����	fF��A�n�a���Iۤ�0�)+<ʾL 6�^��l]TA/Q�eF��MJ����'��䩩�1g6V���>wPm�M�wYl ���Ϧ�,s���A��g��I���A[���6�A��~��IE��X�;i���+�oOg{�w�l>������X4�����O���hn0i�Ķ�5������]����r�����V˪M7�j�>��o���X���?�a�>(�����g�myT>��{��ID���p\Ia�c��v�N�,�F���hX��|쏾�T�<�)[~A��Fi���mC��,6l���vX/*1鍟���r��+�2	yׇ?*��{d:�ߌ�T5��gd;(�jտ��{��{��|	{YG=�L��|r�)h6m�-�|X���hʛe/O���??.��y�ӗ��A���a�'=P��[Wz��h��Fi���D"���P�Y���?'�#H2�����g��%���˥$�̓Rx��0qbNk����.�f�6!���%
��סַ��oU-4[>��ȩ�.ln��l���G�J5�������F0*�:���OL6�6�A��k-؟�b4NZ7a����L�L��կ�Max(Y���Gf��iړ���Q.0�
F0��61��Dg
�ޜ]G�t�H�/ Na��(Tm`����}�A�3ٿ9T!��6F��=f,Bد��"1�!�W�=�D9/��0Ι�F�M Ԭ�
`̘���~�-4�s��a �)&�E*�hP�m�"k�> #)�����}��W�x|8$u�J�~���m	�{���?�/6M���s A���qԺhW�?�H�")���)��ҫ���MV�Y��������9�/���Ak��������{1(aPl��������{�}�THVE�d5)�&gd�^Pu��5�^(�/���8��cr���0F��{"%�]��p��S�`�+��ŽӬ%+����^�J�i��� ��9�I[`��OX���<p9��b���
U��Rٱk�E�� ͐'�+�?�m9z����>�ɻ�}C��%y�Q��ӛ��>$��J�5GFV�#|�[�7"ly�J����bovV��
����q�&�B��1ćWG1'n3�L�E��p�gm��4l]�����tC9�S!D�!
��;W�S�'�q��;aF�ڬIeuӟ�������G/�ìdص} .��{�\��M���EJ����Ӡ=rpD�]�0+���P'�ek[�,�ը& )!�wt,'h���(�oh�;�o�<�YN�Tx-���h�_��w��y	ɬ��P�Ea.����>[,Ծ��ɬ	ܜ�y���)hsɐ��B��ȋoF�L�2�YV��-�-h͔�¶d�� whlb2��ƺ6ٰ~L`>0Q����� ,��.�i����p�mf�R��fir~*X�)����6��"�.�ڇ��So�$�k�H˞/J�T�4�`��0����7ˁ�a��S��A9s����#6��� ��﫺]6����Z0��F^P��g.Hk���=%뺣���'�-%�8O�q`�&^h�kYS=e��J�w���i�f/j�7�*&��$�-�8hJK��:��'�A��'?(_�ʿ���<sI����n'��	L�o�%��5{P4�^lo��i�����mk�L�sfN ���v�y��<�w��������?��ˍʘm�iW���㆝�My�=�ב�,o�F�d�8������=ٻ�A�0�
O��C���� C�rˎF	Bːo~���}�씜�F�E:<[c�sӪ��5�T����:j��8��DQ��TKg�W��`3���G�g��k���fE�
h.;���)P�$G@�=��H?�%����?��!g
�'�E�֟���,����,O� m��\8&���,�j�@�ٻe\�; }�ߒ�'�A;Am1��
x�i�lj��e�0�fX���<�����}I��<+��#��ן�מ�y��(��-��Y2$��
���w��)7�j�G{^.\�/_TM�Uu��5LT5����,����t�{��C���r��G��㸭2���"�%��r]�2�j�M�/� N�9S�K����+﹬=P���ŊY��DABQj]��7K;��CFu
���B\��j9p��hh閎�;��uijm�h�7�i����Z\j�ߊ���)$��m�&!x�Z�&�v�>@P��?��|��B�OacE��Ht����Q�er�тS%�`^���ۣ�g�f��N�H&���f"Iy�Ҵ���rA�y�w�.�֯�	E�TƆMp��	^�%-D�}L�J'U��SIۇ)o8�-�
 1�K�lr��/6`r�T�����8��d�0}<_��;ASh��q> ~��#Ԅ�?�R��LG��1�=�@�-�k��XgD^�S�ı����Dm���4B;���%��u?�)����22��Q��+�Y�g�C��� 4Q��֟�q�������뚙�&ʇB��l,�q2Q������rVy�xPb�q��yP���b������ny�;vI�7���}���� �!�[3�l��N�M�D?H&��i�f���T���yZuǻ5���qV�uȰqi���[��a\6m]-�o�$�x@���;Kϲ�+��i���#+=P���1�#�^��fJa�*>
�#�(���[e��(¯Gez�o�gz:�څc4
�����mm����䧇��0'8�����|}�n�����w��bCb��oE lu���t�$ :��WON�7��U�8A�:�[|54����x��X#;���	q�h����fY��	�N�xW�����䥰���" N8����aLOܸ	S�L�����*`��}�A"���a��G'��؀nsH�S�ﱜ�KA�|��v���#�Q��	a�K�1��Jk�x�z��B�������9	C��q�A	�9���2��Y�b�b�_�+^����u-�I��R��F?506Y'��^�于ײQ5��H4F�;
%�@8��uv
A1���h$P"P� ���{�q�N�4�Sh�&#�ԴP��z�UR���Y5��.V�������M��/�ȵ�O����K�j��4��rF�c=��oC�@=����f:9��.Y��-�aHz�)��.�9}�W0!Ǉ�d�{������b�,���S��^�8g���B�y-t�J����IhZ�9$��iK7A)y�v*����ȅ�H���(
Q�r5��S5�Iuc�k|��υeb'��%
@=q9�?���ڞfTͤ���?��o�ţRW�(�M�;�S���
���KMF��T��A2i6�i��^��;7�ͷ�|y�S-�N��S'�ɶ��I@bn�w
f
ڲ��!n�7��  @�4oѨ��h.q>��T� G��.���9kb\K��gFr9M5���pT�EBAij�x����e��Ǽ��I�i��Ma?�!�x=�Q .�I��0�����N�����-'���A�'gݦ@�c�0�Ģ���1|r��t�1ƥ����H͒�d��U^	�	���d��<�C��;66`�����i^��Ot�,|���:&�o���	17fF��a��Z!��:�χ�џ���I���UmH��L�B 85΢@��chx��4���D-�1�)�gj*�6s'8,����0�(q�j��^尢o��v���|���]�e�fH�92���4.k|AimƻZ�˭��'C� ^�P�CY@9�u!�]�x�s�ؗf��$����^��~9���xܸ���AZU4��"-ЪpU�i���m3\ȍ��	c��4R���籪vx�vJ������:��j�
B�'s-���_���"�}Y��KOˉ#o�N��Hg.���?4�����x"!��[���o���>_���yRn�J�����M&���̼��i�)~;�YB�u����&'dj��4�dϮ� $�'�s!�'�B��[� ��[ev��ׯ��[ץ�D���8,g��:"DL*���~��� ���['.ȹ�ܹI���(B�����G�W�m��vL�c���O��|O�����hv��9؟ r)��cIR���Ĩ��]ݪZg���<.ky	5�j�C��(���%��l��m7ɛsd�����7��[��NN�I����2-��wԍ@����s�b�/f�c	��ji�M�yղ�)���L�0�Q#�9C%j��U��	8x��>��&�K�D�BU� �Lmt&O����E�`�����Qߣ2vuK�̛,�:uh'���ݰ0/5j�٣�u��p�|�>�g�X_�3>���4#ݭ"��)8���ӷ�6�@�D��PЃ��^�J�
���jq�>gn�V�����ȟ�Iy�'/�zߜ�b�%(IH��=Ai��mLʅ���e�yɊs#�]|i�����Ѝ���j;O��v���Ɯ`�5QZz�j،3wA���HFb��c��@y��@���5��j���ƻ�,���ܴ�Q~�K������'�;#��<�($��!��!��Gv��޷��&�߇��gޒ�y�W���&��K�i��o�{�5��&-jP���[�ċ��A���yZ�|����ʉg���>4q�/��(��	h��!h�J�2[Z�t��S5EhX���f0  
1��4�,%aZvj3�zU�_��S'nh��K�a�_>z�N������o�[���r�G��4oy���r�wF�MO�l��Al�6[�~֎��_����aÏ����C�0і��̤J`:�i�34��9��a���&>�Igy!�����9_l��f&�%�{2J�q��bj�,�CPg9�;Q#5\�=��)��]�w ����.
a�b��N�!G��G����"�;#V50ň�M�G�A���R�k�L���}���Vܧ�Ѝ����y;CE��H�����̕����iΏ������W��`Gvd��V������X�
\����r�57+r\�Gc����G�q1���&*����B']��y��y��@�]:�235!�C����Ba~�-����䣛V�Q���H��汷�F�S��M�;�q�\xt�6lJG��!��v����1�l���['�|nF޺8��zi��ͩ��O�����LH�N퉲LC��f�ذ��t?�r���#��S�m����I���[�/��l%:��Mù���E�n�c�%�����E����-T?���Mr�����W�i..�K�v�ܝ[�\[��꫇��~� 84����޺�/����Pn�9�l�+�B��d���L37`%�)�*C��#����Z,h��'��B��a�>͐�֐%��)Ε:�8�8X�3���ay��<�T̹��BZ��.�GM�Pg�	�x�1�fT���vJ�mB?��2���+=�ֆ*i���*��C�4K�W
��҂�3��J�\w�b�0�����e�yE�TFg]��E�ѹ�a|VI�5bRX�=��h��-�Z!U_]C������ؾ_ $�&`��Pr�E�:��q�&)n�����C�R�F??.AZ��p��5#bV��M�H~b����>��}f:.cL�N�%�0̨�8��SMeu2}���<F9��f�j`��~�}��tX��`�U ���::�8����P�b0�K��j�XgI@K�e�-R��~Ra�ggsTe��}��W��'}���r�>U�pM�Q�l?�	�/�R�߹�k�
�C���9A���9F��,KJ�hbZ�՞k�	sCy �*����ƆQ~e3Mn�9��,͌Q��w
����\N TahRI樁��J��N��4�K�a�6��b�?m..����D�Ւ�m��x���%%�ĥ1���1��e�L��n�������Ƞ���W&�?*c�pI(1��X:��@���0Qj3/saP&P�鶐F���Ne#C�\}Պ��eo]�q�v�'��NlZ\��h��֟�D1?����\bjn-$�����%�3������'ic����y�e�V7w&'���MM#y�<��f8����.�=��顡�Y��w�Ϝs�ڜ9�D������LozC�6�)/���.�z>� �t�61�qӫ�Ɩu0�ԹŪ=�f:27�y���<86�fH|Zʫ?�<677����`�1��l���nt�&E�!�m#u��̡o�>�Բ��#�:�7"�״!L��N�\�SPQ��W��0�L�K�S3$�IXO��p0�3�����hs�d�ī� �	3@�{������sXk�dМŹJ`L-��s��$"d��21���V�S���
����#C��}P~0«��)��^�}���fIM\������ODo�T#����Sy���tlWS��J��Z�Q�Ҫ潏�]Hl����y��A�I�Z=-��{pX٦\m�����` A�'#!�Q��3��Z�2ƹQI��/z9�b9"ŀR�7�`�~�
`Ź{�>���F�p��U��f���?�9�ij��"5[��\�p�0+e
����:��Wئ���Z�3\��^�1Q���"Q&}jy3Q��|�k�����L_nD6�b�1y��s}r�"6hK�q�&Rhy��]W�M���׻�h�K��C���7��\�4��Ŏ]�������<��Mkd2*�>y��ʅMj�A{���͛��&�JU���'&�o�ڱ�����1D9�xld��͘�G���2�v8��9�(=���e�o����Jn�dӮC�S}q�tL��/�����KH4���r#�(��iDO�K4yM���cG=���n:󗞽�qa�:?#����� S��g��t'hin�33��K]��;����Y��\���� '������%[6���u�s��d�j�>݃sA$l�ghHP0@˔'��Tu�{�G�}�s�2��X_��ۺ��������<'g�\�]����>���_�/8�c-(�?A�V���k�C������b/��ߴ�N��v�O8	�^�S���aZ݂54z�J>�ul���}XZ��2S�^���!��ۈM�f�NW����\,�<~��u���Kg���t��Z�j�<�j��
���Dpf^Σ��v\���S.��h^�G�75�M; De�i;�;:S-A�Ei@�U�{�,w%�4�z�4K�LX974�Ĭ~'�Q-�9���rss�<x�;��V�����J��81s�^�n��c�{AQ�A�X���L����۳[z`ɢy��P�a�kHӐ6W�C���&����G@ GF�i�|��K�({�q5CO��ASwk�z��( �L$V�$7O�Ͽ9�(�1i`��oN�f�"I�?�����1���;3��`B���7������4�14��e�FA���U����:��Վܷ��|`<.-�qfFw�������{��8>�vx^H�u�ļK`�v���]��偻����a���k_�^=#��ye���@��V�^���,n�PW�*t�.'c����k���h����]7B>��O��]��?��?�Sǎ˖��KϮ��@�S�sP���F��L�F����#���0W�V9@<5!��9��{����_b�!]�P
���9:���)cB�9��	9���B�v�</k�fĻ�+�R��X)K�+&�����l5�\���g(=�FA��f��� ��W�:,�y�x6Z����N�D�/���r�rJ-�H�q��A�1P��q8�s3!�N>-[��ưm�.�Y�� ��Ƨ�#菉tS�W��A��u���a��˛�hF�9�^���*MM�ҦN��!	L�I_�o�Y	u�1�諊Ŏ�fvX6�J9O1�ي?�M�����	h�Md��*2"�;�@9��0W��ބ�~|7�Cjr��È�(�rq�.�E����j�Bk܋u��&�by� o!�6��&}�����+緹�@���z�eo'0r�466ȧ?�Y��������!9��)��C���v i'4�.ưV�La;������M����}���cE�њ�.>������_�|l@�ᚂ��o�
[��9L�H�ޙ�mb0�4��|�����Z�Z�`@�������͐��"������+����[}�&�·�	�<5���>.�o>'��Q�-�ĩٲ��d���4�z+W-�V4L�k�V�X�X���}H,VX�s� ���ǐ����-���u�H��l�pD�<�)��<r*� {҄y��)�u��#�\�7��=�<��>�_H�<'���I �eV���6lJ��m��
�xi/�;� 0�kfx���Al[d=6!�T��B����I-H��.70���XZ&��i��5���O~[S���х�ƀ1���Y�� �X�c�6�2�p~�%�QS7U�S(��s�1[+}Y�9[T����?���������Ss��ګ*�RkDl�� a-�{�P�-4�6N������"�e�I%��}�TȾ�#:y��E�5u`�#;������O&8?3��,�8�7imT�dV�u0�����5=�h�b�����4�rm�N9��K���������u��"lm�|�{�|���Y�Ώ�Vy�z�=��ar�Q��e�;�����<�ʴb �&|^�co�$�o9�K>��_7
N�~��U�s#t���	Κ�y.����qf!��%�V��x��A;;��ls}�N26#���c@Y�`����z�u�MU�P9
7p�\=���G���C��!���aR�]�|�9�s#�lˎy�8��,w~��{77I��^.M�F'�>EvL�Q������G3%�[�K9h��zSؘ���
c����^k4�+d4���X�~�#��{��Bw��^�$�T���/�tSb��mn��������S�'a΄326rj2�q�wm�X
9�4_�aⶋ�s�e �������(=>�w�����t�S�� �y�XL���ܪ�ދ�������k+�,�{d�,������ڊ����Udk�܊>'KI�h�����k 2'���m��Z���<��
�O��}r()�7��d�4���M��dn�5ݶ`�b=��aZ��{ &k���MI���m0Ŝs%�#LwI8�Kȶ��s=�� �Nh�j)��T�i�<5�͌�;�\���&>W���i�';��nև�'N#�� ao��&�+ցjB`�-
}r/��)!�VF9$�}ʞ�1����ـԼ3o@2�a_i�kk�x:&`�
I�pV��}�6�n�����!���/��ݐTӆ�ڿ�A�����J�_Gɭ��U}��M]��`@��2��|��ϺZk��Z��^M��6����.-�|�Okd���썙iA\� u�[��!aj�l5��<��R �F'���;��/;ֵH��"}�����������2 f:LZ�Z�s���˯R�׵Ft�ԁ���hJN�p�9#���('�:)�yǃ��[�(c�Q�������)��u ,�a�y��s/��p���
~Fm��!��-p�9uH|m��O�-	��!3� ��tv�%��֯�˯|�l�1�� 2}#Q�����1�$�3����zh�T���Pa�єy!�Jv��_�|LzVI_��.�SI��+����]�r&�c"�lX��\L�0�l]4 ���I34e���7G䚦-���/H��N�Q�8//�i����� '���1��BO&� x��>D�e63h<~��mP�p�|m6P429#�ϜM;�S;3�#�r3Y��@���/�����5��r:	h4��p�eQ�d�w�K�������%�#
��_�鄹����{�\���Z�=7,n`Gk�i�S˙[]X�]gWS��c%�㳭�M�R'L3��l�y��t��y5��)D�oC���i^~�r�I�n�4�v4����"I��+�����$S��j4"�-�ّv�'�P9�X赜vJ��S+G��>;"��6%a��U��*4�u N�����!�$�3�0ߡ/n��&�z 0^� 5rd�~��a978�k�	�7�A
s5G������g�������M��W2�o���1��������s~��Q���P��|G)���;3YJ��N\4��R��r1�]K�^��X1ɹ�k�"��8R;P`������r8Z��rt}�y���$�) &�N�t�[v>x��g�䷿wI��G�*���=Y�5Y��ph�`�;�"Ne4�����˦�7˖M�`N��S����
!�'����ɜB��P[���.����!��:�j8su=��ݏ|lkH�� ���k��5�m���ldF�R3��e�GƝ'�u�M%%[�n�;n�%KBԕ�4�������H�i�dר��Z~�>#x�}fӴ���� ���U�}�h7.�~��?�����3j�q΍��vy�"��b�^D�iJ*G���OZj�j~��`}�W�����Hl�(R�`��Q����"?8b�I�j�HyP�dS�+� ��6��=6k�&���I`���!���ϩQ)$L��~������<nw�n��w�(R�BM���rv D�&-��CS��ѝ�C�8����y$j9R;�/U�yKp��߅�ٗ��+���v���ieJ��̛��r�����l������K�f��@����g�92��v��D�U��[WG7����S�~6lB�����Y'�����#�r&ѧ)�u�p�#b���8	��XEL�=��;v�;n�A��[5� �֚444�c7��ȷt�M�������A ��n4�6A��XJ�)�fGh�Y��fFs@S�3峗ؑ�w�6n(���]w�����MfY	�,���n�Zٷ�z���F���Ry�o<���FG�mTq���2� bժ6�����������k���u:,�C��,9s�U\��o��4+���Q��
$uB�c_ ��h�
��M��� T��\|�7E5�����B�Y�^����0O��5e�1�k��@��C�H��F��Be����r� �ky�ݶ]�ٌ�AZ��	ծ31�Y�r�O9��-�����1�ٷ;�.�'/U[��m͎�uB�.(8���_%AS��u=���p텆���Ip�D5)�,~(Ы���w��C��"���/�qQ"S�z�7� �}�m��26���H2�kb&-�0ʡ���@-}���Z��ak�b��l��7M�8�)uD��
�Ml��t���.^]��qx� �����J62d��{� L��!�G�.�a����]��1�U�)�9���t��v�`�F��(�&'����e���"�F�Qd�|Z�\b�R�X��F~� ��ƚ��8YR����5R$�LYBM0�Gdj��j"���\��gAت��H����ɊAF�"��<�Lk �?Yf�MeS�8�+�*�+��������W�sB�^J�V�P �^��c����%�S��Y���t�i����K�䥶��{�F#P��A�7Ġ�7	6�$ԜW[��ՐoK@����L��"�L��s����z �3� +��Y�<��)|�q3�F�ƹ5%��s�U�<;��A��@��Z��M�z���kZd�َLJ���N�D��D&F2�s��ln��Fn�5xg�gBHNƪ憅����9ÂΒ����"���j&���CH%���	��t�p"�(=���s ௃&u��E��P�|K'�P�~7	�+�?��jj_\�&�/ ������.���$z�gw��ߤ�1~a����O�L$�#G/J�=��GIt�����;R��ޕ��s���Q�5�Q�vF%GGy��B��|@��Ƥ�u������>4��ou�ǓHR�)`FGz���	�#j�W�r�kB�TeEô��*�Æi���EXR�3 ��$�/��Bߕԛ���0�8��ԋU����)�=^�nm�b�3aCX�S���(n6`�&	��ؒ��Y
4�%����+��=
A�ҝ�^���3��t��m�A�����	�!�U
��֪�(�^�%���d+:8L�868 æ�]�*�����<uu���y]A�&>��95{������$S��fi��U�'A�`�k������ �:0_�6m�³�N��ZV0H�Ĕ5��_�|��86nچy�9ݑ�V��r�ʳƶ�Z��\�999�j�U���I�c�F]�߭>a�[����Ӥ���#r��s��O}X��{d�m5��Ѯ=B+����I��:�Ⱦ�u����}����鈛�33 pA ��^�����.�����>)����to�\�{�K)���}�9+cç1O�r�ɉ�VM�ť������̈́k�Iy�e\�4��f�Z��f���k��)�2 �'�⥟�h\--�Ɲ�Cd����?�1�k�H�x��\%�?���`
Br$��"�;[��k2�>J�(μx����#�u0?�gg��(���å/����h���;%�Hy2�k�Ԟ<����A��|?�E�O9�FƑ*�,ָ�����O�_)��g�	�1��N�VF��z�� �J�P�{L45�[,s�Ꞟ�����4�~:��9ʜ��>�_��<�C9��"3�[��^e�""j�Ԥ��KK�0�p,G���D���)�[��-uQ�qо����4��|V`�D>�\�y�Q�^��i�h9��j��'Ӄ�khz�߬yY�z�Y��o[�|�I����W~	�4[5�K�,@����J�����ʹ���$'�$g���Ⅿ#�f�����9�u��B9[�Dٌ����R��d/�i�\�XL�����UA`v�j��N�Y�|*Zx��c�z�l>��I�#���&���6'����n\θ�.BY�u/MALIA`���'un���/�Ǎc��*��g��9vaR�,�kHSH0�MN���xH��<%��P�&3�dY���x��K��_ah�}
�� �'��,��I_do���~0AZ-AZ6l"� �+�2�5䩰�x��+�1f���Hi�����V)�j�'���� +���A�5�m���k�~��OMS�uRJ���� ��!$�U:�R��m�s��A$�UT�,z�E�en��uhhPN�:_(j7�y�X���j�an����-5��n��Dȫ/�����QY��qI5��C겅 �g##2}�i%	ݼy�̵�$�3�΢'X^���V=�� ��۰.A{(<�����ĸ�I`�]F�$����!-� g�(^�����	Q�,2:M�\�5^�H9�-����H7%�����]L�P@n�h�|@���tʼM7��7@0w0!��WS�&G�a��{�������KGO�l��La�pv�0̊1�o�շ�sC3��Y2s-����Lk�w<�ci�Gn
�b����o
����i�3���A>��/�a$ZΧ���2Ա�5��f�w��q��;��8����a[7N���Z�+�i�mM�,�(�@FV}�D�T�Q�B�*�o���)�r�q�܌Y�k�hR稳�꣄_h��o�&? �e�`��'�2��74�S��o~�ǚV%�,SF[� z#�����!����SJs�Ғ��C��>� �p(��A�K�zfZ�G�9�*��3�
h�Z���n��-M��/Ü�~oP>|۬<|>�p���Z�!����?J^�Z{�g>-�5?m��ί���0���K_��7,��	B!� 7@�PazMXв4�����<ǚ~�����5��3M
Bz��~��y��*:�����V�l�^歚K^5f,*�t'��:�o�|R���|3B�����JA MV� ̃����輻�3dzNЋŝ�*�&?��AM�y@���,�aJ�0s:�	�2_�'
�>�;��w�}���CG?+�4k��A��.
�����I9�n��P�S&Z���?���p ��������V'x�ؕ�~9q���EfX����̬�ߜC��48N����8##?B��y��F�k�6��I���P�JMLIM��>�{	^o��ː~r�ڇ:�ӷ+M��|���΢<p�Z���+DD�'O�3�)�����`ھ>"Uu�C��w���f�v�3A��Q�I���:�\��{܃�F��D�Q�"`ڞM�1� ,r��������O.I��I����6�ʻ>�>	6����=��a9~�On:p�y�{25=Mݬ<�ċ��ǫZ ���/����)�JK�k�wV�m�9H���~�a�F|�}���&򲌁�ЙB�	�tS�	��n3�t'U�$2	SxӇ`�@= Iӄ������B�5��_xp�l�3�S3�r��9�-'�H$
b�� @�γ�r�Z�����ݱ^�G���#nHC�k ���[���D� ��8���ȷ���)|�RS�=���r��K3�����2�@n�d���̥�CQ9v~FMAy|���SS�`sc��a�B7���
��Y�?<��� ���sp+�����׈iJ�JuȖSǐ��Y�����4��H�R����R�K����\�<\0 ���Z�#8(̹)mp=���+G�d�w~x����-)�9Qäf�E,�!��#9n�@�2��!��vH`c�v+^�Q����22����R�w�U�R��/�_�(�4����"�5v�,��Zr�::�fB�}�{� �~�cp��%S�a]���z~���� `bZ���MA�|���������,OXL�-���'c4��s��$��?��-M���`5U:E4Zn���kUK���N���[d��m�*���_�ǿ.�}�B( �c�x��<��������@8������{x���Y�?���B�~�M�q��ǣJ�&ᐹ�rޘ�v�q�3�.W�aoLn7�B5�M��X ���T�V�BzD��Ƭɰq}b.���me4�o �[�C�q�V��Hm�2_A��B�ߐ�Nמ3w ���uRwPq�}�69�Í�:��c����(R�*�R��+�f��2}!��Ë8\�ٳW�|�I9v�����#y�Ǐ�|2ua�9�L&�Ļ���o�W���� ao�J�k���)�j=��X4���V.�ÛW6m]#w��A9j�L�Jd�R\����W&�Wh\u��E4�M�M��?|V�@v�%l
H�ʓ�17=�dҦ���{���u�T�c��2���o	iQp�2�. �;�"�%{՟�L�z*��x��i�<0#ã89#�C��=b�(@-�&H�
7�쐎��j��/c={e�\��2�Z�,K���T�l��1�r�qΫY�%���Z|Ov�g��y"��P�p�#]>�6�h��S/*�6䙚.~r~���ϔ�	�B�禰6���Z���_ejt�Q��ʹ�)��š������~|dP�3��ϵx�
�i5#�l7%�������R���ɵAX��>���5z��Mrn��۰V��h�
V��_3���>L�!Ҙ�� �Ue�e��<O��8
P��#%So}C�>����O�}�M� �΂? ����S���/�##5g� ��&{cM?����lG��r��@`�c��Aa�2</��TN�V�U؊�D�,<�?��\D�]���<0�U��e�bF+�����S����9j)�1�r� 1����e.@򐱰~d��^\�?���ƮE�\�܇�r���4�m5��s�U�ϙ�N�J9�i�n8��MM��3�/�o��\X��U���;����OZ��7ߣ.38X���[��U�*����+y{� 7�Z� Y�Q.�B!�l=�0�Y�a�}��Oc�p?�5z��Iy���&7�|�> ����g�Ʌ~��q� �J�Aa�Sp�� �Cs��	�P��B�� �b�{+U���x��F����M滃CHM$5 ��1z|J�$7l$��f�
9��ma�@rѹW#ǲ
4��f�y���o�>yp��Q��\t[{�-��v_�1"�&��~�"�k`�Z� �i���	���Ji+P�PY�ʃ���T��T�C��3�s�Y�X:��cZ7W�_�>rۗ��M�!������W��G��\�U��JW9���]�qۇo�� �=��,�ܦ,cc�_�m¦���Y��Eqg�j�	��I/����;��g��%9�T7S~�_���������_[VIc�06�IM�I� �[�5�n�$�'#İ)9�U0�nέ�cm���P`.�*���[h��F��:�I�n��{�-j*I�HSY��SC�QW��K��s�U�#��p�+U?���E� R8��\�=&��A���������CQu�^�i�hR��s2JM�#�In{L��3�&5��@���FJMP
��d�n�>C9��?v�Z��3��c��+�~��-�;剳�rr�������j5�h�ZZf�m�����!��٠�_�z�	�K͆�߫�#��'��y�{�G�y�4y�;�����L(�E���4�0l�B������ܾS��YN�&:=Y��aU���PT%C24�/��o��#|���T�����Y�N00,�C��pu̵ޒ���/
V������Uz)n�L���i]-FY�
6����/FW�5��F��L�P�}N��{c����)��'$޶KB���h�jS��V������Lr>�^�,Wâ��gĺ�dѫ~?�Ч�X��`�(Q�o��=' ��%�}�rh�f���Pj��O0�g�U�:�j�.M`���j�r5 �Oj@?��P'��Г�l���֢P2i�ԁZ4;�R��:* �l��U<�Vn\F=�[�����O����n�,K˨�+UY=@ �����0�ղ~s�l�[%�� �DA�^L|b�^��q@v�[�����C��i�^���י�^���'RZ��� �y��6%��&�BbU�B����X2��o��9탢�1:n�Y�č���%�w��jx�=-�!*�ܼ��	�f�b^=�c�p���}.7� 4��� \��*�T+U��G
*�� E@%��o����=����]
أy���ߐ��O�\�D{�
^������m����~����!���N3�:�Ҽ%`���fk=4MQ������l�
�M� ����r�_��1 ��ȳ�8�����=��H2Q0}�x[	�K�$�屈��Y��,��zh�%\Xx4���?��_	|O�3��1��`TeU�EE��%�!< ��_P��)����]�'9��O�|7�$�H���k������:���&\���$��j"@^S<lf"�-����H��z��ɚ�Q���ȿ�ӷ@�fLq3��8��0A���P-�#��O���ٻGn��Gt�K'�;?�,@�k�*L\�g+3�����⹳h���Y�0�,��^��ۅ���>5B�~�P���FH�?�}�,џ�&3n�)h����A�r� ̙��{7��B_5Т��N�{6�ʍ�o�&\/c3a�ޡ�����6L��1f=�
�Xݖ��߂��@��I�;��s�����'ߔW���m��M�0X�e��-�r4I)p�||��&� ���52��Z	���\�ľ��}�8jJe	D���N��],Z}��7�S�9�нI�ٶe���w#�_]�.ª�F�"V�偵rz8OF�Jٹ&��-s��5�m�e&�>}�� `��	�{������gU���QLʜܢkɻa�lJ��:8��Vo��I��=�|��e���z6�e�(��+�_m=@�(H+#���}��@a�>�k��yJ���v�����X&<�7٩ �����s�q����Q&�-PDc�r���)#������r�m�ȩ��<���w�+
�t?�"��}��|(�M*��ϝ;ki�����/��/kt̷~֏\kH�A�VG�u����p��I4&�=y��d��[!�A�	%-���7�L��� ۹
�R=���� XjFBԚ�((�V>��3��(�(7c�ɻ)��igN޷cD��ݲv�V�5���}S�8� ؔ�f����0�jCx~�x���PP:@m��QƦ�2n%s��a�{�>Sv��ĉL���#5��=���w�m�+�����گ���p0�!'~~�
K/�3�2Ce��k'�`����c�D�J�zE���2�8�]���/~B��9�Lgi�,D̥?�SC�eJm'�0��]v�?�lr�uc���c�?"����'�=���[��qٽ��rv��V~��Y.�v��r�3����,�
u�Vo��2煊���(���m}���iA
|���DH^x�_9�x2-T���]����q�p*|j#��:MfS42�B�f"j���aD�ٳg��u {�݂M�	u)��d�(�?�M� B�Pr��4R��L7��j��<g����R݄4־������#�/�@��d��X'�=�u'!�LȰ:��c3��l��N�ע�>j���S���ᔻ%pH���C����nh��r���\Fz�/'�OJ�VpL	$��uҳfC��Z��u��i�<��+h?��j���� ��9�?-k:;�����(r&v��`ꢯ�b���6�k�s����i46��|��#:s�-��F���tw�8��[�Ɗ}r��Landx��i��� h��oh�&s��k�Z�)�y�F5�ơ7���>}Hb:�-d:��a��ʊ�͘>��%��P��tGq��_���q�(Cq�5˼錤�G�;<���˓��_�E�G�I�嗶v��ԍ�R��\w�1��6���\�/�HM��O�&��1s����U�=b0-���>O �P1���$�����q����ՙ�Eto��k��(HҦ��&�M9� ��aesG��6���r��yh��o���q���K�;�P"��^=�u�<QG�x3/��s#	�)�m0����Vy�����
#�u�[@j��{l3��X�&!cg^������|���uG��fJN����ȱO��J9js|i
 \� p���$4.6 M��y�(���2��'�K#�r�oQ��
�c��ܤ�۠��3�_��~p�fbV�+�-��/s�!��2��;:�'k�`�w%i��/�F���];�M�I`��&�L�A;KRV��`l|�sF��b���5E@��=���� Im����a���w���|����A5��������&-�l��C�,xH c ��W�6��$��!�?^��|ڪ�:��];������[�C��dd�2s�˳ߜ����zD�"��xćt;L��n+� �7�����!���˸�e��]�ރ*xƊ���N�o!AO5(&�<8�	�S�hz��<��9�a�c�*&���}T�2�H�YQ�Xߥ�?U�k�Mw|���ȏ\��݃��؄�i���1��lP��
��.j��c`����,i��s�.�&r��b��L�7�̆`Kjj��t @�UurH�§dǶd����E�3rÖNy孠� ��/{�a��L�g��nج��t6ť�1)'�c��Ѡj?8�aWbWP�!��Њdm��\��pr�D�[*y#��~�Ɇ�0�,O��LD�d,ڬ�� �0d��6�8 *�闻�.h荦�fl�� @�:����Kr��#�c����.Qԍ$�!pA�B�O�:iF�&����jd�Ŭ;l�ؙh���^�ߡ�J���vj���H�����0��T�:�P�B��"h
��r���F�"�W3��<��p=�ƚ����5��`�~�c��L�U�%�e���K��t�j��W��8�,����7�kF�?5ʫg��z[�%W~_�w� Q�����6ET��i&"ra4!�B����0��G�.�C�ۧ�X#�pg�*F�Q�8'6�[$�[��޷C~�fH�G�h.*���n��J%k�m�S�`ݠ���h�B��ɚ�3��<*4	����{����W���pV��C��f/��g�}������!n��vT��^h,��n�f��LP�*���cC���T<!�!40	��sj�J>��l蘋qe4W|?4}��چO�������ͱ|BM5����;:��-���g�yR���_J��/b�����L|��RV3/����5�n�X�u|�1aW˖��|��n��4��ߖ7�-���\.ŷ�_���p��6��Pi��g-6�_�E�"�,K��U�(��"�
+�ZQ�3���y���]U�hK���@
^F�2Y��ܙm��䇇����Y����t=��|@�G��D� G��Oj=�=!_�ޟ��D��"��='ݷ}���ʟ�5�ڽi0]�c_^���	�h�W�K�?j��
�t5}E#�s�v��L@ Дa@�
$�)���9FX��>:��kR0!!�wU�M Ҋ��5H�Q3���;(U!�T�?��ɏ���tƤ�Te����rM�l�e���K-}~b8��Uߩ� ga��u>$��L��m��e�Ŏ�c�c*Y-�̼_6�H0����-ښ:�O5�Ul��o�8���N� 5��#���)'�I��[VwIK{;~D���5��o=!�>i��C`F��o�tX}[�Rk\9�\�R�0��ɗ��?��}��}�i�~7�J���/��0�AN�5�ϫ.�!��z�!�m�qS�l�~�[��NP�{ʻ�9���9��މ�z���T�Sծ��?yprr����Fh��%����I������~�j��Tu����p[��O���{��#Һ/(���Cg-���u�5v5�]�V4L���W�\��<�B�D l�X�A�'&&����&kG}�%���s��p�e\\����(�Z#���_�L8
Ҿl���t�!��,�⫐Nf�j�ș���X�A8��S��{�lݺӪ&�6.?=4)��55D�	��r0��0�r���~��EW}�����]om�������Z!��<0�ܲa��y�pXA�I[^[8_S���N��y�$�+cN�j�"]Dj
>/,��d���Oay�w�*c=�]��	n����F��0��jo5G "Y'@q9AZ�*>��.�3��S9�b����U�v�q<�	�}"�#x��� �w���0��p
�`F�gwu7�yd������쯴�t#��D������x����f`���8>g�S�(ɍ�/�LA��]�P,|K>���M(�'���JC#Sr��V6\�(a�9|.,g�S�7U���EX9�$4�[��f|.95,��E�ng�>���3G�>�I��j
ք�j*\��������4ψ�]:/�����Ўy��ʒ�]���̀>���}�o�zy�g��% ;�\/�t��Z��C����&�hiZ���v��Ed42���p�&��b�~x�|�����j�p��l��d��6R;M�+qg����hJK`�Ġ	�qa�7�9�אƢ�����	���:ٺ��ʠ]����J��B�˾׍�v1�s���b%�������wH�޳Gx�D�GvsDqV��vF��7Jզ��W�x�+��I�@��Y$�}�G���5���֥�������'L��k�ޣ�	��;�rC`%ӁI-m4*�����#/"�>t�[޹�[�����;)�����F��k��s�	�Ю��Q���/!�OHl���N\�Pǻ������y��+�XWةK��tc����ف���k����l��I�a7�g�D���~f�W���8\�?7�<�gحR�c�e�\�H�Hx
?���q�3_��/.�i�z�ϡ��_Lt�F�p�zm�lڶ9Kf��@���g\�o��G�U�Z�0�J�P9�ZG�w����+Y?3�9	�o`�c�¯����D}.B�|DF������In)��m�lj���?�������!׎L,��9wR�ly�u���r9�.Ǯf�07'��Sk�8O�Ŵ ����9��(E���
�Q��G�s�ps�1�Ttϳ�L�JM@2R�	��d|�n��`��o����[�a�k�N�t����^���Q�!�A��>O4����_>3,��IS�e
L��0]&�q������B�25�	�E`扂0��7��װM��"e�<�ǥ~1�F���0�)!� )��l9m)�ZR�N�#H��Y�\
ܡ7ɋ/>/����ey�{�U_�(= ��J��S�O��V���˓ǒ��X�֊f_��B��)SfS52Y�Qj|3C)h��Go�v*��,e�t�����)́b^Y��[�Ay;=�����_s^��Y���P*���"�C�l0�j���|��r�8f�/���sw�2�a2<-LQU�d�z5��1/nF��U�T�L��Aec��I BS#i�c���>� �
�?��f��q�t0�Ɂ,�tv�3��L`3I�G�|@�����D2�Wf�.�R��:\�My~"&�7�6k��&�l�,�|n�;�c�x��%a�I���E ����PN/W�n黀o��	S�1��G�W��|�5h;Y���~��=1K ��`�]��]��P#TM�j�
A#�����z��l���*�#�U�P���#$i��s�ȯ�d.9��+�G6��[��u�˙�#C�{�zeQ^C�Y��X�l]��8�yXh�h�������3�����X�5(9L�i`c-
a���F�\,LL�Q�Pmύ�6�#�",u���t�^�$�֋Ӣ+�E��Y[W���F�:��9 �$�Vf=��P*�B�7�fa����R���sEb�y+�����h��Ⱦ��q6n��8�	P��^�*s �ī<��ω>K4M =��d���˟�Tt�"���x��ܽ<I��� �ghSM&"�6A�^����;[��W���taba� �<R�9�h�c�ܑl�&���D�M�����j����pc�aD��)^{�"wG��#ͷ�r��Y�nj�4ҶD��Inѡ�\���	�s�KQ� 9�Y��C��򭟆���T]����Bա:^.�2pW]1+��]g]�Wq{�+�("�����CKb�ZX|d,�IP
hT�Ä��֋��T��h&DZџ�m
 e�0a�\{�dR��l�T�'�S��4v�	M�����l�O�7�����#�\�2'�(���R�-�S���-.+~�d��qY�.*�?�[�f�}�r����=2UkĒ��aH|�%�Z,M�j��.�WNS�/�`�&�=r6&�p/�Q{��M ��(";2��3*�D���n��8���$�E��U��%lr�e,�k�u�8O���ч˼9Z���Ls+�3��Ń������ۻ�t�P��^�X�/H������ȅ��	�$�惈_�-Wi;V�[�XL�חo�'a���kZ�{@�V��ؐ<�mY��k�E�]�2���NV�YDy�P2/h�P�)+�O��ouO�1QqS0t.�7b���#c2y�GH�4y'��΍7�PӔ[�ü;��v�+}�	d�#j�i��. �LMVi���3�:^�G�I Ǒ`֍����Q|3*��k �$p��J!�ԡ�����M��D�a��t��Ⱥv�##ri	s1W#`O搄�P9�6����\su�@ת.پ�_�>��0��a2+�Y��e�Y�d�Lmj�I���s�4#9�^��׆�����J��Ȩ�^�"��2p澺GpQk����Oߞ3ĕ�oj�F4��� ������U6n	ˡ'|��A��2{�^Fiqc���B?�ǥf8�[ё�ͦL3��Ҍ���DyVT_�=� Z���k21tZ&��4�VIǃEju��z���J}5�q S�Cr��|_R`i�����*�ʜ]va�eG~=M_�5�H��y�h�Lt\e��ϕ:1����v�dЂ!.����O��������'�����ʟ|�kr^nB{�¿f�<m�Ī�_!������گ:_�4��ﲿ��3�7�%�<��T�ۮ��ϡ�¿qp9ߡ�����y ��Qw�!�o�� �C�9ˬ�YE�%QRU�A��K��]�~}.@���{.w�Ze�aAw�s�����s�;T�!*mb�*�♣i��k����\��VZ�ܵ�� h`8X��5$�4>I�0�n�i���j �U���r���
`Z��|�>���<-&�F!����H�u�|�d�0MU���DX�O�:#�7�,Ղc|?�Fq�.ٶ�.c��洌g�52��{�d�8���)psȗB�k�������!�nB�[����9@��JQB��r^N���Ah����ɭ�ȿ��-pl�1�΂?i��l�F�D�'w�9�4��1���zqZw�s�iSQa��[��)	M&sx�Ͱ �v1�/lkH�;w������,M��e�u�����j�+@��<7,|���M���D��j�0b#��˹����&Dn_ۈ��9�h�9��KC �3<�mj�M��5I���蜼plD&��<�V<c��V$�#)�п��C���i]�:륫5�\A^$f;gfr�줌�.l�-�����T�N���H/d�V����h���V�c��Dߴji�����xF�	�g����c�
4�Ĝ�hrTx����(�����sn̕���TpV���Ƴ�E�I+��a ���/��oIS�N�o ��{�Uw#x���N�\a�Vn��V��*�k�..t

&�NX<=�̄���Pk��5{:	���ĕ��N�559>���vlh�w��d��y���L.��RKe|6 �<f婟 ���v����,�\w������ d�f��?�e+��,�~����1� L, X�.o_� �S�H&H6}K��a��r��Ϣ�P��S���!VSE㿠b��<9&A0��m��Gg���s5�e�j {�����h����e�
�wԾ���	S���'�ɋ����<!�����w����� �h+���^�o��t�q���Vy�M�
�X��8�;)c 5�(� �>zw��0��^=���	➤�[�;v���;���1S����22�Q>�:���!����0��)0h�\߀z�X��,ܳr������E�ի) N�E��
�����r�����\�:Ԉ#Ȃ�a X�@I0��4�U���[>w�R+�6���8SG�?���V��F��R.g�h�.go_���!G��뮃�^I,�$���������g�T�_����H����-��(8:�jd[��-uFZ��|3�`vi<����G�oH֯_+�m�@�EJ��*i������lٲZ�y� 6�����v/�!C���1�_����+�K ��h������L3���Ș<xH6m� ��z�464��s�>����}��w��ϖ3�he�m�A7�¤�43�݇vPy���7!��+!  ��7(CD6mUʆ,pn0�-�Z�jlg�];D��jx�������9=��ơ���`����@O�'���(�F�����m4�tX���44�p�`p�&��L�vO��bC���ŶƐ2>�b�(�Qo��UK�`����]+�-�p2������u�X���ʇ�	�=U��*Ǚ|N��K���"�M�+ڨ��dw��YLe�ص|)��4X��84 �G���(ξ����oj�T�p���-~h�#����V0��4\�8&��ۮ~�TU#_[5ѳ� �?;�ӧޒ��Q��&�w)%�M�qɼ�-�]wބ����oG��kf�O�ٔ׭_#۶nTb>�M��1V�i8�db|XΝ=����1d��x�vp^].*=�"�6��17�Fn��"�La��\�ʣ� j����>��X��͠�HHd:�ה��ȁ��Rdf�F����� �A��R���B�,h��s�=ׂ�=�L|}.��G
fr��!VH��վ�YIj�	��,��|?b�`�c�z���g��c�;9�S��E���Z�o�OU��p��`Z��a��k?���Q�CJ��w~V��{eZ�<��Z��\�V ���p�<$����7^�ɴ+���~���#1�
p���PK�U�3	*�obH;A�7SU��|c�[	5!�O}<�Wq:-�Z;:ז��î����3�C����d��&��}�9���V�J&tu�� κs�E#�-�s�L�#������z�b��Ѐ�[�{Z�R�Uz%5A��<�V� �o�=W�Q@C��L���~��٪_ɪ-�v��ݵU����]���բ�f�m_���%5�^�ܻ�F��?,���X���N%d���^����%�����\Fb�׃��u����ǉ�~�k�����σ�pBpl��;��k��1��箅��:�p0��P2D��S��6�j��ɯ��IWN�����B#iS��u0���5~9A��P8��>\j�"� ѾUGǌ,�Ga������%�M��&;��H�j�f ���.�6�Ś���Ь-U����-�+A��r��꿥���E��I�J�����G�>gpfA'���IQ�:{��
��Y���/w�!���Ôۣ��S�>T���U�����l���&� 0qJ���d�۹z��E����
`*�ۮ��S@G��*�w[�Z�ޱ6N=�8B�M��ɅK��U-}�Fu����W���ͨ�κ O)��l�2ޜ��S�}�]��횘
��?O�v�@�Vb)��B��ӈ���W��J�
l21�FQ{d�D�Z���C��"+�p�5Z�lJ�ӑL��rR�ע��\چ�=���� S�t��$K$ihuu��3ߛg�58 ����|Rs��gd{qM�
��UW��2�d��z�4c����|��c����ܘ�,h�׮j�s�_V���0�d}�q�Kp�L�g��|�(��Z�Ս���M?�4��Ü��,p�0��5�Iǰ�I�i�����^�T�9�Zn�������t�ܢnS+����
�ߎ�N�N�XlJ����4�J>-p�f:����c���+�$	���cH���ʰknh<�FQ�k����Y�����g�M�QR7��ͯ��]�k�������4��d�(I�����=���4�9�ʉ͓�M{����T�P��QS�Vs��&���N� 2lGj{L�e��<&����l����� 6�a A�`�`0���`{Vf�jh�P��ĵ�J!��� ��P�,�ʿ���Q8\{k�����uF��D���h��D��9�F�!�]5��<hl��,�<�}ҍ�g~��:0��L��8�����v��f�Ĩ;�@Q�l�C�Bd��M�����O�NP�O�a63+v�k��G�j��J�}��.)��@#m],���ķ�$փQ��V,T'�wp2.�훧�=��:P>��E�� ���������h4�������j^-[��_%{���T�q �X�]t��%��;�Z���i.��ol���p�]b8o��,�z���X�L^BFI��M"Q�CpFRMBa��G����߼��/̉?],[���ֶV� t> ����wJ5<-p�i~||Z��l.�x�?���A�Z�1zdd|J�'fL6�&���7xh� ��7 �O_�M7��]����ؤj��5![�n�uk7���|�t����°!0?��"���f{9B�ki���h�F�l[�Ye����峳���L��\3�6ݶ��Ls24�+����f)M���hJ~��Lc~���l�R=3������Z91�g��G�6ᕦ:È^psai����y�g�����䩺�44��k�[�:�Ip)q�$� h'"�q]�8�)>���� ��Q�<�J�`5Lw$B|�4�2��W����vm���/ӑ*9L���q2,�����ꑠ�>�0�9+Ӄ���(����3+�ꐬ�ZEO6�تe�Ts�J���z\9��ؤ`n�3;*�3?�R�E�y �<�Nb�� �<P�;:�3`���J15^N-�+#��x�,|&ə0��&2WMZ��&R�a�8	#0�	�x�:�;d���]�a*�L a����'-��D=�e�w\�+Qr�E��ΰ�.K__�/Q�=87��MRpଊDbz��������2�58ssX0;:�?T �\� @?�\Фl�T�S��9^V1|���l�!�n �9Ѩa�I�K,��56�(���������ҋนE]q�.R�����r�ޭ�)DI�3�g/��Q�"��B���,4?�ޣ��5˿����3�h����m��Ϝ���*]�oQG�6�a�ŗ����;�cd"��L!�G�I���*�QT�qY�"�+��$�H���{l�_���;�>�#͜����vp��p���o�7m;���B���K��#��]I\� @&|�{q�7�_��1��%�:�y?{�1�ߙ���(['� J�y&��#U9���3�䤒��(��9d���� �:�|�ׂq�ț�~�F�	�&�;a��I9����_��Ve�������P��F�kh�V���hY*	�|A+~�G��#�䝖S�/IH$W�[-�A�,����d�g��& ���v0��͘e�ђ���5g����0�j~Ʊ�]�l3n���z�C�Q{�[lQf�������
�)Z�)}1 X�sF�����
>�憺\�B�Y1�]����^�~8OOMɾn�֖��5�,r^��e��W�Fb�� � L�r�Y��2M��f�]��}Lk!IaIg\U��A�Jz��r�\м��>��clvQ�s�LhN�<�;�T�4�70&���R0XʌD�v��-��{�i]�(?r��~�.��y��#2<:yՌ1�$�������0��1��F�����0sku���Ơ���@'|;�~�;ʮ#�mGk+o��\����)Z%��ve�@�yF�$@���e:��������E6kE�ww��&�<��=��I�˩T����T���%��=P��E牢����	`9W(#��ղu}����?��_�=�w�'�����[%��NF��L$%�9t����#�q��	���'DO�,Z ���:���s �՘�W�-�ރ�B-|.�QM��c�흌X8��@r	PV��
�I{u�O�&T���&ϵj�]�;���+��0
WC���g�I@�T�-F��D�e�S��>��`v����UU�v�w���'Hb�$�_5O����x�U�	B��3�rr��#L����#�IP 2�7j
�,����8L.&�5�
} �h�UzR�&H��lmO��x�V�p��|	ߙ�B�<gԏ��o��Ƒq�^���I�&���ܰP˼�ڑ�d �3�<�����X¦UV�ep�}�[�\@S*醮Zy�>��I�-{o���S�?~��d͝_�����cJ�G����'���=�e�&#@N���1�q�z��沁��N�%4m i��9?C6C�J�a
�Ш��v	� �U3[�d��ګ��,���:�m�b�1�~��N�7�;����S��N%B�C��ɘ_� H��<_~��isO�ɶ�k"Q|�c8ĥe�C�^ �(�K���ɘ��E������j���%g��,7��O�z�_��z��_i�.ٹu]����G ���$�5�q瘼��)�\��g��(|2f�/�ԅ@�T�WR���;h/G�c�����0OALz�96�!3�-R[_&�*�Ԋ�����0�o��Q����]��ji�"��v@^z�5y�C�?~�W���^ֻi>�5�v�'�~3��� �hr�&*O�0P�(��,�78.��.�/�#����}�O���ҧ���>����q�����r����*�i����t=��z(Q%'��GT�q⦚�iț�)�wR
$�K�Pvxav��_��G�Ti�F�z���p���H�n��3.�켄&�+h-( �Þ�
���&�-|�#p�ho�m�{�f��n�hB����^Vu�����s�:���W��60�v5s�7��9���ηO�2�<�Q-@,L�ңͣ���ã�Ia�m_)���^�	?)�a*=��5��	y�g�;���-r"��8廬%5�̑�����w�RP�?��m�!z�c�� ��*��M���u��P�2�ᜟ��q��ݫe.�)?����dD����r�^0ͧ�M�q���;V.��V S�}w��	�l���g�&�|Q��3#�C;C�=C�Z�8!"��Av $:x3$��9X���BfO7�Z'�$^�?{��u�` LGo[��줖��H�SŖ,GqI�?vzb�qb'N��q���[Ͷ(�*$%6�b�%�����;S��߹�ͼ�o l�;��}������/i S �R..�ZRWi{�.,Tˤp�=KX�) ��+Q0��2��(��l�&���D#����A��X���i1�!���)��lo���̯	̅f�*dF&YE	,i9�˅��t��
�)����ezc�]G�<�6�!#�X��ߕX����K`�n9;ڄ��ٴ���0p��[d׆ZdL�e��0��I9xfD�	�&��+�^0sy���9*OWP�u�&d$��t�R�CXC����?����]]S��* ���P]�)qU2��2��xL`�������-M�G�Z%�D��WC�9@H���[�`k}��wK�1L��86�$�Ĝh��UJլr�+1�Cu�H.r̔shjwA�9�)\Zjԍ�]���2��VVh�g�.pX9�rE�-wrEZT����0E�Qp��¼���Rn@:7�W���� �VA�@�A����<�@�U�������q����A�~�VU��!+@ũ�ot��9TΥu��z��Y��E��,o��� (���2��:w��
Z�%�r�&u�%1�W^���b}Oˆ���}׿���~�#�)�������-y��d��-��/Kv4M�BN(�k|>�U��'�	�ώ�jw�݂a��hX��-��/���[j` ���=7 �1Ѣ�0I'`1�5+C2��Sm��ܞ$�+Y�Rc���S �*����+��s��ȩ�H�����z�YpƲ6!�#�?8zE�[��^�g�c���L�04�8����� D��lgK��>�x��H�(R�,��58�L�ÌH U���Sܽ��XW�n/*b��$28���*,��`Jb����tߍMRB�o���;i��ֶQ[��3	�,�I��l�|Vl�M��X�	����������֝V���+�]j
��5[%C��Ԅ�Ie�N����O7�$o�7���r�)�z2"�oIo߀45�n��j�����ij]�w���TDj����Y|ܵ��`)nfP"!e	�z�x1[�1��6m_ 5� �<U� �4.�|���M�Z�uRy6����E �� ���{���M�^�T ,��������3r�b_^��=}��ЙU"��s�����am{P	-�FB���a��P�ǂ`ncdG&O�������]� ZM]�wN�M:�~���\�L�`�IeQ��`8 ]�J,kÿ�+�d]�+?q�ry`W��Ɖ�k x.vv�_�ٟ�޴<~���A���0��si�
�Z`�,�
"����`ٟ>�%+Ο���[d�\|�)����(�o	ޡ	 �B1�j��#�f�����>�hm�Tנs��j�Ż1<,_������]Rx��������.�;]�xI*Ah�l[�.}Z�%|��[_���B�G
��[6���'����!�X�R�K�`��a
/�4�O���\*4��Ҕ���ޕϘ���-R7���}'�9.7�� � ��@�S�=q�S��;&��੗2m�Ҏ��uw�]*�dNW�O��.�S��ܚ��Յb��	�嗠���|ą�V�\��r=�Js��:y��e���k�T`+����L��<;�H2��Ke�V4�8wa�Dw*�����{��};S��j�G56:&�g_��G>���d���iK���w����q5 (G�������z�@9��ߔ���*ڲc��wl����|�]ڧ$<�'/>��\<{Jv��a�n~̸�<p�r!�kZĠ�|qTJ���l\тsaqC?M��/�&�w|%��V�rc� ���E�܂鹿$���0@O�`��Ŗ�z�~s8���3 �,���m��2y	�^�1{AA�9�#��4�qZ��</�N]���0�Chځ���o���4�ٮ��'���,�[���:��wy�g�.Λ�BL�] Mu��4`�2@�@c���AJeS��x&3�� lQ�Y�qό��]��K�<c͏HrǦ:�cKXvnh�����Pp��/���$\[-?��Yw!��������d �E�'��>�@����c/��.�A�;Ys�����E�;VI��Cf@[b����[W���f��׾ G���_�?����݋K��N�����;�w�&����C-Kڐ��-SY��/�)��y_��}�� 5���Iy�.d Q�{�!�)>�GL�ܦ��z� ��,s�)KV�9h����6��FM�3Y{�`T�7��Ng?Ǚf-;�p	FxM��D�Ȍ��ftY��������26�4�Ch5u���!���BW:ZXj��{aˑۗ��_�쓝��T0�ʇ ������?'ǎ�����
`)��6�L��;{ޓ����x��J�x��aL�e��t]cN� �$��q��lڤs7��O3Ȱ#xѹ�7e�p(,M<;`��@�u5��C�����	c�FgP��`��P�R��}GɘH��+��r��Y� h��`� ������:]����o�"?5��c38�x��tr8��_v-(���>���|���gj\�M٘>4�7%�	r ���5k�����[m�SJZ������p�Bn]߬�7�z[��1�DM�0FD�Km+��9_bj�����MƪD��zrύhy��=�9�u����
l�D���� c��ݍ��v/��2�j3��7�cFmF�:>�a�<r[+2uk���/��oɑ#���?&��m���#�Ա��S�����o�x�T��K*P��I[H�?�!��wiʲr7\��=��Qy�{/��G�=<>y�@ �R�ae�=�6'��e���t��ý\#�۴������jւ<y��{A{�K����A��E����j	��������M�o�%E�Z�(x�FQ|�+j�R1�<�Z�;�塛����̓u����Uj�Σj)������}ظͻږ���R�}<��T�z�m��V�K7Yc�&k�O��?��`׊� ʉF���BI�3�ݐ��l"�������(��O��L��.�q�Hȹ�(��;�İ��mkD�=���C��r�,��#$�$e|)�ʋ���n���X��������M�73Ovb��D���#��йQd>N��~h�|��+��C��#�<��A�BQ�'�xR�;��jMG.H`���]���IL�|��L��4�µ �UTX8P&�|xD�N���}�,	����_N6�q�̶o�e8�����I�-��1��rx���m[�u��w��g�8�=
)���r��1�/X��I�	�ҧ��t=ԃ��D�bv���ņ�@D�Z�Zo�vɔ�LN&L9�/2-����x[�_���&	!na���R_Wg,M� �}�܄��)9p�Z�L���q�=�ڽ��������` �Ѱ��=2�%��d�:���ɳ�q�Zٵs���a�C��x硰�em��q��)�M�͂<�� Ufk��eɚ��@����ԛ���\�;266�ҽ]�>/��1���Xqy�{zL�ǻ0�0�\�;��I.kųeo�#����vk%�-��zfR,A{O�H�zd�-w"�혼�����[���A��_��_��L�-WM�D�O#�H��C�<�w��(�c`}�Q�� ��߃�&�]�a�qه$�OX#�TQ~��:)L���+��s}2�"�v_�g�Y��ū��.��i�< L�PP�"CFh���,��������훚  r��+
JhU�v4�nꔟ�1J 8<^������>h��r̼KZQ�5�jì��Z�����O>&۶������)}�Ú�����v ��G��C��͘NOűa$%�i^M��[j�|�֬FaԀ�x�b��7л�-������rcƜca���]¸3G��'�]���M����f��޵�8 ^#`3�п\�����^�5�RD狑���^���M0�,Y�s�,t�E�-�/���}�2sC�|��?-gO��|���o��g1�	8��� �r�T�����Y���"�n�(ʪASRҕ�x(��,����Oh�`ݲ�2�.?���b�˩?�[��T �.�=�t�k����!Q���Cm�����@�6��R���iű]5��l@5�;�15��+я��U�?��� ��m�q�BKK���w�����1��w��窆��sE�H7`�����=A2K��Hdh����7�����_��ԅ���. ��iF=8��q��dY�unYI6�%��������	�̋e^��(���6�S�c��}�2Y���'�c�j��מ �,x��R.�im�;�_&��=;;���[�d��&��8��P��� �`��<��'�o|W^���O���h��
g��I��w���z��V�i���a�pd�md��
c�T ���X���h�?�ה��*ʛ��\<r{@y��mY��*F�$�D`.7�_J�$����g�Z�>�#f6�Xw�E��oKǢ&?��@�@�6�=��C	�Q�_���.y�Ѐ1҅�rI�>��!0'qd,�\�� K�~����n���$Zs�+�s62��o��)'/F�[�����ץc)b-����h��;�s�e��%ds�Mr��J�z��E�%�)r5��sL"k����r����# $�x�_���4����(�Ř�qsZ��&�Far�9���r�����\K�*~��X�W�sMxANKS������� ���Ȉ��F���Mf`by`��'���]CƼ̍�J�>x.�����]� ��ޢo��J&m�DK ���h�&w���e�r;&�L	G��	z�SY��"��������-�b##��R���UU�|���ˋ��R[%� Nc(�͹BQ���ƅ@#�D�`co�,K��3!���%C
jI�5Y�լ阎j���Z�q������j�����{r����Z+�
�3ٔ}�����ʽ�m���f��S�r��s�o
���@��u�?pn���]��Әs1uFY�'9�1Nłf ���/���qY��C^�K� ���c��v�}\��B�G��WV�Q���{�:��I%?;~�2��)��t�Xj����P���/�v�2}Ss%h�+�2S�5
�g܇��4���n�H�T<��d����|��v/�� w��N�j���)ո	�&��L#f�g�\�7Vw�e�*s�4!�
㦩AЮa�<`,L0���d�� ��~��r~���+�]��D	�I�Z"��e�&���gW����:/�T58_�<�����8���M�N�x���֨[u�O���;��[_���NY�tI���Id|>����s?�9 "��M���C���!yq���鼧�j7�;Ѣ�� ;�ዕr칧��t�ʎr�C����p6��z��79�-�|��tKcs�l��Qjߏ�r��������7��`�y�������ٶ� ���r@��z��`J?,�4���=��_��2� e� jm}�k��(��-;P�"��
1�Ȝ�Q�|j#Z��~�!5�5�@QM1�TZ@�uqT��@>y������z�RE��^X ���R����{ ���E�di�2Y�t%6�F @�t%�%`���[2c1�ÖD�5�鳛At!�P�0 H��8\,+��H��x<����ײ(	g9p���E��V$0g7gʓ$dd0"a�Ju��e��
� q�l���
5��A
]b�H��e�S�kU9�`]����y�N ��2���������ܤw����>��p�x�\ʗ�ڰ��c���(o� m����MhP�S���f��INvNɲ�>/��v3��Y�q��[�,�d^�H P-�n�{_�Cz��D�:����,�p�f"�?M����6�6�e�(��s�p���/���$�D����2�|����
 � ��f��1V�b�VF.�G�-V��(�Y~���-/cl�(h��KKcZ�t�9!�#lG�mtd����~eA����ݻ�-���!������-�d�Ͳ�����z��L#F�}��tm�cvq�K���X+�|^���'A�G�?gƕZ��215�9�e�������M�҃zg�;4��+�`�7�e;kȱ�	��kX�4%��*e���2��6{�#X"�$�Qg��(�,�s�T,������i ��J]cX�{�^��_����)���k;��<���/���2&��6�r�{�z�T+����,g��#�	�{Uk��c����xZ]�W[LWz���|_�3rw['���D�ƦT��s���1�Vv�OɾH�đ�9;�AC�I9����)�J��Zr�li�Y5��J�Xj��!Z*�~�/d�?�@�Zp4]z��u�/�e�{��|�?��һ �b��7�F	�O��\/R�TNTʹ���/1���B��\&��6I�76���|�\@���Z�%c�-$�F�j���ٲ��	��QL��xzo���sE�m��x�5��^p21ƌ4  ڱIp����5�h����J��X����k+cw�ǉ�H2ָ���?-G�w^yI6m\'��ܧd��5Xb�]����K���蹈��3��`}�ZY	��9f��o��@�_���E>�W�>,��#�6��[��^BHd  \<.K,������C����}Y�4.�;��#dF�LV��6ӝ7����r�\3��`���VJs4�G�R�Z5 �K��ɞ��9�G���V�Q����n��TN˩�Z���R��n�g��gF����f�8��R[��z��d3:E7���=���%vfO{�� u�8J�g'�Ob��D���kx��a�}�{�l��u;;f�bq �J����Ҋ]��q�	��V�iV'�&�)2w���d���3 FW-��Ѹ5eۉ Sc�2,U�m���	­�����O��2`�M7��\��j
.ڙ�P᫐�闿{�h)��������;��1~��c�T�A̍�+ջ���F�;�����'����uȠ���q���Ku�||�H�0�� �am��h�H�E3F�#��T-��a��_!�{���h�������!�	%�:���ФN��`έ�jV-��/�۳R7�l�t5���P��0�H!�͊.�f�(����L�bv'6�)X�"��m��"h��5TKs;��-�L��;�l[�(?,KK���(9�!g?X-E��&�g���3���Jd�&/���X3�iٓ�s��4��wz�V�O��?�g~�]�������q.� ,(����c#��=�N��U����Ʃ�f	��/>%_���'����{n���}24ݘ*�2�e�M8\'��?	[�e=ҟ�"���E�\���ki���Sii�c4����+�f=��0�-��@�d|���BMY=�y��A01��U�:�`�"m��-w���@F&�����Z��g��{�~��nZ��  cA���ب�]b ���O�fQ^�sM5��az��z�}W��Ω���_���9yn_���2��I(�)�{�a!�.��:Pr&��ٖ%Z�	WC���8=	�.��:*��$���ԛH���:��_���/��:z^n�i�T�b�����=}C�wS�cl�	I�e_ܾ5,�H�E��}���ɽ���+%���*{b��n��ٝ5������'>����]������ɧi]6�r�,i��N��y!��b�
o���z7��V�i��%�a*+�	S�&�5�K���S�`×�.�2�f\K��=�#]"L����C�[�4� ��n�L` � ������A����<{N/}}_\N����&���i�!H�@E�cF�P�M��-Ct�f�^;e�Cg�� r2�J����9Dw[�3�#>�����'����<I!�Z��}�v��aXŪ��Y�M#��Am����(�5�t"Y����W��ڬ�ӘA�s�"fж�+��5�`%Z�
u]�9G���%���<�R���n�Yd�N/�K1"��=����W���vl8��3=�9w���?%�0������� P�����ik��}�îZ|�Y���s�P\߉�������6B���g��8R��|��T��.l����Adb�ͦ�r݈�3z�4>D� a|�G��[��6�P�9�����,0e��i�,��5N��$bt���Zh�f���S`��<;*{���7��O܏8M|��[����A9=�.�+|Fů����+'�c�^Wo����d|<"��~Y��U벬�x�Eכr��qY��C:֬��������Z����Q�_��=f}&��4����rA�"`�u�/�Y�r02-�}_�e@~�{�v�xr�$ȑ�����Jo5e6��z���mA��R@�'xb@�q�5�v�i��|�J����`2�Zd��~�y�7��� ��]�$^L!�&�f�ٖ����<�e����KQ�=e�%�,�%�,`dd49�2q�sn�IrE�"�����[����pA�A��C[8G��3�[�1o�����j^/7��>i]�J��N9Y'��V��W�E��-�r��!y�&���e`�jy��&o�l p+Di��	#P;���bdb;���.m{���2_�a���ji�&��uɑ�a����vlH��-2p�Tg/⥫eX��vPp���y��r��3�J�
rԒ� ������ �h�+�����/�>}�x�^�֢ζ��l�8P\b R�6{����4"Y�Bٵ��HpLy��_}� o��),�ˋ�a�ZW�ҫ�F6h�#I���<�����z��³�/��q��j��[$x�ؤOjZ?$����]%�x0��i^�t�S�{SR��ژ޾�gT"�r磇@��Lj�c�eB�=�F�D��i$����]�q� ��-���/Z��O��;r	Ü�{�x���wV�	�� U�
yw�N�(�x,��|�������ϩ�ǰ)>7K�Y.����#c��3�-]X�3<L3H��W:O"�9my��Y�����uP���%�D���8�d�fB	-@��p�}� ���S `�o�*Q���h7�L��`���V;�5+e��O�>���jHT��c&+ [�t����/�����V���A�˗�Ɂ#[(J����LJ�������~����%����S��cW�m홻��Wj���2��;nX)Kڗ��i~UaB]��O;%S���!�ЙC��k���f���?���ե����tK����ס��kh\z�ߝx�`�}ll\I7���fv/c�Y;��j��0��~ϺZ�#�Lò4ɂ�� q���$ My��U:�{nl�ma��|M�����\F+�o���Jp* W+?�-�t3�wDZ�a�a �m�� �0��
�2C3�ZLO��9�ue��}`�n]�$��!�0��;7���2¯���.J�~�m�ɓ�{BΞ<-�M>i|J���/l�����t�f�ha�f���6T��X�QII��TE�&��� ���}I�\<rz^m�[�$8����*��gx�x��P�� y��83�_����(��,�:`�q���pk������i�� ؔ1r�>*�LЙ�O������f��zւ�����>0�5}K�c��9���ٮ��/ɳ4� Kt�q�Y�x=�ǒJ�۶D6�h��Fv�;o���e����\���`n�*ONV�k�<M��i�<%�R5�B��jD�۱��y�[6���Ѝ��-�zoS�%��C�A�wvJdd��O�aA
\#�庡# _�:'C=e^����ʮ�M���J���/��[$���]|�<�i��8v��?~�`�5�U$2&�6n�B�s=(,���� ӵs_լ�iZ�Lzx �
Of>�NS�u0��G
D\��J^��� 6����ZM�DB��f�ϧ�F�Nt�h�v��iM��ƌ��$b9����԰���![����� `�dhi���̈����T�kqn�λr��)�����fd19�=�N�$GD��q���V�b��eCP�gx�P�q�qG"����c"S��	J�#�i�Y��$�O�%���;2~�va��EJP:::,�pc���~�*u�&�y9Qh2��l�W� W�\`R�)	�9��mu�l���[��+�yB.zY����G�V0�O�����R�̴Ip�R�	n�eN��%#���{��C��P�ߢ ����Z��q9z`��t9z�zx� ��m3(sRh�j�0�e2���G/�t����"�ܔ
��L=݄���OS�;�`�$)����~� � ���X%�`�����@��e">�Byb4��G���t�o�@|�C�f���@
�8���I�E�j��-���(��0���l`1X���3�1$`b�K 4�)��<��/����j�[��!V�	�P�plPz�#��_0v&���sza���ׅ���d<�¶f�I��Yy�̈x��@i��UK�:L��8�5-�����O�0H�%E��
K�M��'�и���]�U+��M?*���$2�X�LE�Y%�!O�_�,�<��ذ;݅y\)�����Ç�y�}�B���No
Bs=��9e:w<����� h.�s�WjX�Q*#R���>(Su��"����l�b�=��\v��iF�SA��	�nL6r���o�=��p�J���d�h]�J�J_��������F镱HL¨@~��]r�;R��S�
� �hT��q]�sB���*�^Ox��k�L�tк3���{ޔ�����Ȑ���ɮ�[e˦��cm�80 '��^�ea�&`)��)VZ��U��D��4��%, Id�M 0M����X�*l�~��Ț��#@����~�X"+���i�@�ep���v��5?.�X.7�0M �*�-Ob���k2���bu��� �r�\��ѷ>�/�R�<�A�CPE���T;��x�C���26b�e@�^=�d�^��o�3c��r�g䕗_�#O�Xg��%�>�ɗ���>�s�\Pt��s>ۇZݴoLg�W�o��}^. ؇C>�[�M��Y0/��.�0/�{�\r�v��C��|i{@�(�� �(H)ti!rU=W������������ �U\���]r��qini§�9[(�����Ɔ����;�(���ɍ��o�w�*��gL�k��q��A���eKBpg!&�s�N��ưQT��H@A�ssa�3���mWi�;�0���r㜄[�
.9u� ��.����ɺ\i����>���� ��`s 0��0�	"��+-�K��DP���jI& �\�t�:���9Z���B��6����	�`�$��=S ;�'<�S�`�*�5y�6�R� ��Y�|��Sr�GjCuR��e���ڭ��i��Rb�s�N���d���@��F{�)e�Mm`�W�1[f�cV�(J�y��%��QR,�.���J+����-L�����.�q���j���m�iܯ,�L!��eú�(��!��R0w�̀��G�/7�����Io�4���p͟L��z�
�㎝�2�7�T1����Z��!$A�Wz{�@�͗�C �K�@�n�4��#�M�ma .]pA�� @d �V��`���t%{@'��m��&�#s3��5�Y�v��~�p��I�����&���%��˱��$�w� �����:s;��}��՘#�&�R�✌�������M(9��AK���D����qY��A�sӄ퐮�̨�i���*�c �u�G
 �˔�H��������k �i���J`���X�0�.�+� -Z�.�H\��i��)�*̰*౻$oob��;�9�5XY5��>��z���Sg2��ڨ�yIx���F��D��T�ة�V&�0%�� ��sƩQkΝ�c�N���7EN��@C�Q�Kl$u�
u�8"ſ��.ye�Pj��s M��r�)��/�X�y�����w�x�8\M�T7���:Ta�xQ��X��3� α��S��O�0��.����$�]��0�w.���°RU���}�߄��|�C���4X2�ʼ�G&;׼��/%����j��(T"snr�"�����⵮z`��䪛O�p�D&Ȧ����N]W���}����%u�����(]-t?ekr��5�]�.#( ʫ�C���v��$���yF�$��89����@p��5���1X,x9xG�qe��R%w�ؔ�#�xjf8�ki��ã� O0p�z��~��(@��a�<M0�Zw�$���0�,�l�7��k��+�b�Ǧ%^ٵ.���Յ՝�:�`j�H^��w^�Rw�:�	��F��|*���i��,lm�9��Z����Jvm].^��{4����	��k��F0yWT���UH4�r?k���qE{`0]��vN7��ˍu�)�)�J*<Y��/��.9�R�j�7W7=�	&�8�c8�[l��s��s�#Q�;"�R6x�tiK�7 ��:���߫S��Db�7%��q�'��V 8�փ�F��h%�~eӝ6�R�5au#�gx�b������Gjr�c�`խ���4r�ѵ�5��r]��G�X�n�J2ng�^���OG��_C-8f��T�W�\�͉�A���u����JvuB8sn��hkk����Jne��/n�G�@�		yW��e��Ր{�MΘ�uX�3���L�|�}}f<����w��GꛔDjZ� �Ehb	�6�����n�?��(���P��\����ҭ S���j������͵��tOfo,ʴ�$�Us̙QH���lLlH摟u�`飑�Ƴ��F�&�U��qJ΃�K��H�7���!Q"ۖ��:��ҼZ6ҟ�U�P%v�l�������4��3��lPK/io�@z �m��?A 7~��A	��q�Jy��y�MK�"������]r���*��yg��̆��f Q��lÕ���h��,��y�D�:?�O<22��������ִ��*��O�ǶOYשk��2�E�+�R����~��7���9ʼh������b��K�����Ykkd�Z�w�Q���V̐y�����,
\z*�u���u��ɣ���Q���oZ �:WV�t �A���m���z5����2Lk�z�vf�h�o�[x"�~�h4.]��������*F����~'d�-�i�VY�lv�y�
jSn�M.���Ԍ4l.,pj+�������#�7b����5 B~SN��K:ǣV�]?HM�`k�+(8�������㜏ߵD��	+��}��EF��<!��i� �¼�*�g���w�ɏ�F}3	� �/��[~�s��
�n����'] �#�`׹ԭu�s���̬g��tL��r��9��i�_�Eڶ}@Fb5)k�&�ɒ@L���J�[_���Ҹ��P#�PPS!��)���J������$��A���##�W�9Z�͇�RRbh�d����̗�+��*�}2�u��2��1�BnX㑽_�#y��/H(�[�����|F�a\]�Z6o�|�H�)S,���WA�ysd+���.�`�G-�Y?�A���%�`���aFb3��h�wgD(,�F'�$��0@ �$[",�	b׋Đ~[w���a�$�����s��"����0<#_��W䝽�ʅ󝈭����݀Ӳ��ko��o�O��?��ˀ���1��h�Y�>h�a���~98��o��UGr����l#���h�	 �p��Nk\K�ܑ1�B�<��V^@��l���8R_��#�	��Ͳ
�;ˤ�{+ca���neH6�\L<8���DB3�nI66�j+b�����{W����Eei Q���aED�֧,R��n0Ǩ��S+���A ��a���+9���ĘEՈ2�f2�}�������/�K���{�}_�
Kx�C��q��=�Q��ߒ�|��R��|bE����	&&���lo������'�>���������V�]�S�^��̹��

�O>�S'�I}}����5*t�H�z��n��=gj�v��ų����_�7=(O[~Y�x>,��?x������D�X��?�VZ[����ꆗ�K�4�ȝ=pF�Z�2�<}�&�9�/{� -������V�M�w�`�MI)�7���7����3��`��d�8��q9x�O�`����(��kZ�L�����Kt��I܊V%j�5�N��;9i&��M�]s��o�may���0�|5&�)w^V`�2���rC�yq4�ɲZxA�@��y�͚[/]�W�e�1�р^X+8V.�x��|��������>*۷oJ�.��Q���Xw�]l<�c���?\YThm�ħ�ó_&��AԒ�݁��6��ʜt��C�U�	>&G��[V��9� �I��^-��>�����6.�x7u"[>@����r������W����dUǲ�"����\�c�:��L��-���o�<�q��JXT��Z��䚞.W}�)�l���-��W]l�\{��$9wj|a��S2�Bv#nZ��y# ��'f��J$�*gv��t���ҼN��=��,ԃ�� �{��tY��Pj���:k�#�����Ƭ V��E�����m�uAӵ�	q�xhY�کYP�p�_'��:aؼ��c�w��Z�_m�J�DO��)���g��4|�ϭ�6�m�ޔC#AݭgdZ��c٦\�d>��H�[o�*?x��O�W�K��3�1����#U�l�y{��������3�4������?xI����w�p�P�%_���_����'���Lt��{񗱰�SR��ae�9Oz����3W+	ƃ���-�'�8�4:�'�+K�,NW=@��G��	��p1�Ej��D\��ME�o]=�:)c+g?+p�3��˹i9-��ε{#_�\�^Rw�GLǕh��&���A73�H#�̈́�N�'�ͽ�1M����P
��d���5�H�.7��)j�u��������{�ħ�rL����?���QCЎm�0)#��'�c�Rkk�,]�$�2CP6U�L�d' 5�ȴh�y&>+୔g���?zB�/}D���93}���@q�b�ؾ~s>��Y	�$e��:�r�������SI�g��
ƻ����={e������~�]Ҳ�C"Z{єw�����d&����P(�g΃����x��߼�$� 0�qn����}��'r��1��ظ���,׺�v\��Gn�ʂ=@�nj�u1Knq���
�j,����L�V��Z<{���{����0Y)0���Ze�Z\��4��B'0�^󗣃i��@���[���i�q����`}��S�
�$� ��Z�H��8'-�KЄMMِG!K$-gq ��{����9h�|D#� �p={�:î�	1��`�vhH�;
�������-|�
�j�j��Aa;zJ��Ne�Z-%�u�0�JT!>
u1�t��7Dw�=�i�����J����4�/�De�LG������y�i��˽�>w܄4-]-�ϡvbEz�U 3mh�M�ퟐ�?~��{%мNF'���:�u�	 L�`����/]�^%���Sr�Ъ�"�++�}r�L����
���2��Ż�Ӳn�Z�Û���һ9�q]�w��B*������Sj�И g<P�D���H�"�@F��%,XI|�G�!�.9�c���M�=��[v%�0��Ʋs%M��K���1�r��&�雤���h�ap8>c������5;+=\�M�X0c�0�/Ht��k��>��8��H������r&`jhl�'��~��֎�9�U໩��2��'a�1�����B�\�#�F\�,��E�A�M��O�o<��6K%,Qg�iYʵ����X!��U���(0�Rh]b���1��	�]]�)Z��/�2M�j�nƁy<� ��u�_�z\H���`�s3Ӝ��ꬸ�ۍ�J�]ӝ�`O���#&�j�%Զ��LA�|S�&���L1
�yz�|4��Ì���2���5Zk`Q�eiE���J �t[��J�5�O"Kt���7S��<�E{ghn\<����rD��
�H�JȠ{��B��=.��"���I�ӏ�UJ 2��D��Y���i�Ŕ[)~h8���Zɐ���i��_,���p
n
YzH� pg�_�z�<�� 
[�/J������*Eٓ���`�6�"^-�Y���]D��W{fn������r)ޚ���ᜤ+N3�ȱC�d+����W�@p�Pt�U�5�Mn�|�#	+7��������X55>Xr�{&�}�S���]�gp�n�yc��y_Ɛ1L����/�7 ώ���}��jF	ʿ��t�옜9�+Cc�w"Ms�2G�$��<�o��Ҙ��Ĳ�dY ��d2��滑�$�d����I��\~�F靱2��Z�Jɯ��� ��#��68�m�z�y�ލ�1q�MeFc�+��\��u~��B	Yt��>O���盳K�q�S�P!]�۶�2�Y��X��q���
��qV� orؐ�0��f &+BPl5ػ�{Z�
�j�����=�s\Yn�ɉ�����O�?�o�]��b�V�?[V�Cw��*�LG3ҍ��{�%�����E� 3$��=��	6.��hw?�?#X�՞�8��Nz�������4`�i�Y�[��+�	Y�q��>1��/���@D&�����?*(����f�8,��3��9��v�+6��ƃg�=����S�t*�)�s�������ru��i5�b���-bfyI��]�ar���Ewkk��sR��ǧ��H�7'͠�)_3JJ�����+i.�F̒�A�;>��Z.ݿ:��9e5�oP�MP:��0�ifL߰V0�`
 d�ؘv�,9���%�����{�D�Q��nE�+ƗqN�Z�EL��Ape��ɟe�-4%h��r����|8��ٗ�>�flu��?���[�&���ZkZk ۵��P���g�<s���7y$aq-T*���2���}sS�gz�_��
��\n�U����	rR�t���Ec�~�Fijj��HJ���Ȱ��fYb���Ad���T���SҘ^�BN++]�.�{5���l�5wuɣU�;��VA�����,�B �8��Oc�7?�2�rKg��46]0�cc6���Z��5�¦�Pۀ��M���@���1� %A$��̐��5
�i�	i�uH�K V��m������˙%��]�3i�B0�D�폸�����H� ��Cp¹�,�,��d�1X��Z���ըIWJG�,����|`*�d��#�e�B���U�+�V-9�����K���v��~��}�؛��2%]�2<���i�|cA��,�I&&l�)�9>�xj�9��f9<�q���uΜ���됺y��6��Fai�X��� 7�W�j/��{Q�kY����JMV���F6삝�]��L���ց 
,1��J��\�k"�ͳ,�J�V%fL��`�
�QN�J��m��Ɛ�		�����N��{2S�(�|�]��A�J��m���cJa S��$��M�AK7�@A�0����!9J����yv�BԍH\�Z��1��J��=��6L�O�7O੮���(_E~���륹�E�	�P�n���
�'&&AV��-�^y�������d|>�u����NކRB+|���-Q�����9ӝ���=�ƒ_�=.�"������i0[��>��u <U|���T����Ku�l��r^�rNgv���L�;P�A(�S��L���ñ �"	9�����g,@T���A0��M��涵�^6�`X�f ��T�� 8R�n�;Q(2�Y��cGTk������������-W�jN]]��ٟe#���X
�k�Ȱs�RZ�H4`��g	g�ޥi��6��,"=�T��0`���j��zr��浌
� �
�#���ṕ���Z<^|w@#�X3��D́�~%��1p5��@���1��8a�so�Ieʶ��F& ��)�r�	nִV�M˚��oW��F�Y�I�wn��:��A���[�{g; �)�24<,ǏC��1�4H]}�W�����!�OG�﫜�K�d�ƀ�E	���~�-pIA�.k�%K�H��t�ޑ�t�`AK7� <������m�o@�+�g�2>��13C��.t0X*f�67�����5�ÍGq��������阘�o*}�6̹tB�k���\[6�p��.�)�/նY<��g��2{��P��7������*
[B�#c�,GQ	�1]J�t�Ifb�-�s������@Ce!�t҈Y��2 6<4�bv�hd����ϩ��.��fp�X* 9���[CKt#|�{\��YC�wg�Ϛv
z���4�w�	I�FF���I:VX!N�;_���"�illO$k^s>���J=����5��qK �$?�p~�s����qdl�&�U�%�c@le]�?ks%�߄y��u���z��4<6)GϏ ��ǅ@�n1�cO����Ih͉ǐu� H+0���m}r�?�u��(�$�]~$����K�կ}I~�S�U+�RW畿�����_��DHiZ���?=Z#a��;;� ��s���|𱇱j�����o���`�<]G�;�v{ ��QS&�\�=�@+�N-\j�2w46)���u�%��M������#��ꎙi��#���q)���攡��<�݀��8�%S���R��{KN�J�7}I�s����eB�[e��.�����H�m���իC� ���Uʹ�����	���
�7P�K41��S0e�FJ�v��g����ݻO�1���ھm��~��۫����(�y�-7�{��`-3��R.�Kon& ۷l�G>p7��L�T���;���祷�WΜ;'��]�m[7��%a��j��f�u����@�7����
v��rT�[�>��k@/
���Jf�]Z����X'[�p�DE��9U0���2_�?�=^�SW��ʊ��|  M`���ز͈8���)(f1��Λ�[r��5K�Pe�Ē��b���U�i���r�����A1��;6��5
�b0�f��ԁI166.#(�Bw��^֭_+w��fU�(���55(�X%���-/x�X���R���yL�m^��p���J�?�.�A�Y���y{�q��{�]�wg���B>�*�[QI�M��b��^�n���%�9��L��g}N�4�;�\��>EE3���M��ə��Z�܀*%�SPXX[��km����gk�!&et ���ee]��I���Hu�XX&]ה�vn�q!�T�*ls�8������An Z�b�����O���������<�>�׿�_���_S�����x���?�ُaޚX���L�I;b?ƣ+e�����o+�dLD5�%}^VS�\53 �d��B����6�)c���t�sܨ�G�V$����!Y���M�Qb������EƆ�?}��%�2�x̲��X���$xl�Dc�T��w_�g��4.�{N�����ɶ�x1�| ^��땟�G����'O��
�A����N����X�g�Ħ�j��K�[�ӐaV�������l��)��`.��$��h���~�9�����vT$P� F��(��"�?��?'�7���_��i�l�/|똜���@(��l��K�4��[��H@� UU��sV��]�8)�9�%�Uνݢx>�¶�{��/�oC�ڣ��ZU@�V���u>����B\��=$��KGC�,|&�n��FYd�Dߗ��K�#[�f�ڪ�A�G�����p���@�	��s?���%�w���?�l&���j2�5ie�0�˶�(����=��mï���t��5�jU�+d�x��8���P���n���ͤB;/�[\ϰĉ,m��ׇd<b�
�/o�A���Ml!IG��3�e�ۙ���F<N�f�eU�1&�0&����{�)$33�{�|�>���#�T�i͝ ��D&�p��L�SP<�c�+SV��%��7�����4���Dt�U�ڈ3�('@�V��J+�bY��z�5��H/m�˾�ӜKg��F2nf���� ������t��3<��Rӌ��6�IY�.(��e��8-'tJ�ܰt@[�3FAJ�3��ܾ.��Ԝ6&s�W 8�ߑ�0��ê�N��w_'�M�p��EW&�YC�֒䮃��"������ػ���h�2�5���I���!)t׆ųR=`-.����H�#犲�c=��M~Ԉ�ϰ����ޫ!n@��)H�9�$ݫ����fM�&8��-r�fV�X![6oQ��b�<�v@)�d+ 4ߎ\�~�87�`��A�f�YG�V�FX���O�-�e �t\Sɻ�OP� �����>�=�5J���&�O�~uC�7���47g��ZgVFmmU�&�+}�|�`VNJ�a�ԼqD�z����dqvФ�w�$�����8�6?v��W.Iۮ��ҒD�$���a���F霯�d�f�E���98��2���$�X�����ket��vZ�@��*I'@UE7~kqe�)Ƙ�MUL�6�jI���d����|�PC�r�i��X���Q�B"�uk)���3d]��O���\S+�}p~%��eR�[�O�� $���l��lϤ�w��e�F��)��Qܾ���j�RG(B
�B=0����j){�QC-����Kݢ���nZfu�l�C�g�߮����3L�kRc{HN�}P3�"�d�ʕji"�S�YJ��l�}����o�a����ks2�J�ߥ��.7��*�m*��}�ׅ���W�=�%jU26�PO�5~��*br%F.���]hU��B�@d-1`�[�H|ZF+�x̱������	y���&l�z��iJHd�H�QțJ+��X9���E�|U	Xld<Af�hXS���,����J�b�����d{�ɖ�|'��,+kjGsL�)��2!�j��_#�I��e{[=�([��-�y�
ā�n�V���XBV{�����S.�@�F1K�i,L�@`�`��b*�j��d*���;۴b. ��{��v��y�2�̬��\4;Z|uɩ�	)�,,C�q��I64��h5?$9�|D�u�bt�T���̫:���l�(x�ި)�(8+�נ�����zF@��-nr=�9�m���]�Z_&�b��[eE�&̗06/�{z<5~��G��/�x
b��{��a.w�8�t7?�F����P�Q���بǤ6d�������|*E^���.�3</���O�y�,��V���ܢ�� ������%lc�J��U�06R�>W�%2}��00A[Rp9W�8:ܯT��ӫ}u�#^dT����0�d�`�����q.U`4W��`E*%��oQ�T��ϴF��]iY�G�� �@�^�X�.��:c�i��}��_��j�7���N
��ޚ1�|���09�f6�����7͌3J����~Fy���F��/�S)���_�H[���/G��h�	��i�|'u��x<��aL�F=�~������r��Tm���w����4`2�)t	��7J4� b�E�*JkK�q�$��¸�����ի�<���XD�=+-mK5H�Rp��5��p)�p�,X���C���2�1:�5�KB�zs�߃��K��i,�u�=O��i��0��|�K��������9w87&� 龮�   IDAT�,O\��9/mҍ�U6c㱸f���2w�`I�1(PS �:���8��Ws>k��lc()���'� @���I4����,��O:�;>w�x�&�"ır�&����E�'�]ڮv�&�~(,�3� �I�wg��Yր���,�`�U^}�R�T�����ɧ�;��.Q%	�J��DȿT�=����2���sZǆV�R)ɥ7wY�R�@s~�%�z�,����t��߿?�_��X�:)�����eJ����jn��q^Y�B�?�Q��uV[�2g�fkN;.�N�RKS�AN��o�Y~�?�GY�z�Ig&jR�zn��~<.�`A�p���<Q=�H�� ���,ϿY+��0,��"���R�NȆ���ю�6k#�~�	�4�v٢(�aq0������̂S��02I���{�m9��ָ����,��e�D��񎂐26>.���ٰ�!i���m�R�IW����M����ʼ&fh�Z龠�ʹ��-�ai �	�G�#?Ɲ���
��V:�c�;�:o���r���e�y��΃��������;i��d�Z���j��k�lٰR���}���䵷���f���H`��\qG�5��APÔ{��fg��;{�9~~d��[2��Ba�� dK��d���Z���h���]K��]�(�lO� ,��32��~�iAe �0�6�_ 'R(� 3q!3Y�2
7�����3�-*}��</8���a�R�@n��.��?��F�I��^v�s=�]�	�#�����6n���	�S�mmA-L۷o���_��7���n����#�L�����x`��X�&���Bӕu)l�bVA�֍\��ȫ��$��b�`�������B�O
��..��Ll{%J�3��S(,���;Πu�dט�s}��G�( f���+T��^�p�6���1�ՉqX�Fe
��|>���Ք��rT�,���܌�V�x�L�9 ����^t���q� cVc���9�͗@�W�Ȥb���af�yi���AlK#@zL�3d����@q�V����3��u5Υ^�k� bǖUr�-���g��v�(](�}�Lg�B���7���M�,UW;��Cg#r��Hh��`m�F�!c�4��ڀ��� i�xu�Jl7l*7@=����V�10>���Δ6�{8:��R�r��!S��>�u6��7����MSx�5LnnGu�b�1K�*��*F�*�b�pj��,��dN�W% (=|��|�Ԙ/~�RiqkV�~��s�H�t�ù��
���V�/5[�<\/� �wm�f��yE7�"N}U��E�=�6OY�}?
���,�A�o1P��N���A��\,|�
�rn�}��5U&24
#�hu�߭��\O�X��ê�5ȖT�Oɣ�*ʼ��������&?6̇n��d�|�	��e��J����M�y�q�%0 �Ė�l����u�W�xe�_��Q�|$1%�¹?��r�aMH&t36)��$Y#���pn�%��::��LK,3�V�h�%�k�8��s^�6���%ߚ���j�3Z�.,ޛ�p���9�wjX-M�Ȩ�O_{�T�g,��@ed�R�;�e�1&��L$Ue�
,3�E%Ő�lN/�,*& ���l珲ȣ�v��ܙO*C@�9�.��Y�q'PRO�9FpV(.�,񨂥�qT����s��3��N�)9H�'��&�G{{�����a�Y_�.e
J�F�/}��3x�\-/�>u.ϛ���\0��9Bu����6���m�20�BV�˝tW�|�*B�s�@��ʋ7��94�����V������F���K���u]���7��@�dQ�-\|z����ղk�����#�O�7��"��X�>���Zj �� �&FRKո!�ket֌zx�Q}8�9����c�Ju��u�B��dT��y���|� ��C�E�o�
 �O���+w��ad%�TB�s-�= ���-�p�el9��]�������yi�|�f�E�TnO�>�*���?�я�ԏ��T�~(�����n�y��l�#����iז{ͬ��eh�=|'cJ��l3��{-`�W|>pk��U���v>-�wy{@]�%۷ͦ<�_����Q�����6�jPͽ��,�B ��A��$|���-�L��q�]z.�@�o��!݇��$@"X�1���QU]#�jU)��xyG��>�� NK/�A��������ƍ�@��wеҫ���g6ʲ���Q�'G� �e g{k�]f?�Շ.��;�b���b���{\�^��{ �x�w����^zi3&��|Ȼ\��{�0��n�vn���r�7M�l�ۦ��z۬{Ϣ/�y'�iʷ�����ٱ\�;n�A���d����=O�rL둑V*�պX-[���;�����l_��t���B�{�1/}��g�J�s���2�)1T�߼e���ڏd��k���,c�(cS�|�q'�5��;yD�K˒���Ͽ�ǲ�T�t��IR��Ғ�D& �eb���Z������U��wTښje��V�%?�_yWN�u��S��j�-l��3ӭP)���/4�p� ���!y�ʶ�Hw�])Rr@��~SPc�Vhk��VRxv(��{ە$
�k���D�f6�,�=��	�~�W~�G�G��'�x�A��K'w��qP#��t��?W�9�,�.��-�&ż�[�?`&�
��N$��|@�OY�K��p6��_</#OǍ=�����U�?]p0p
f�J*Ľa��m*$� �{�EFFǤ��Q{�Q��n�];w,��,�B`�q@����{q@���|6*���ś���Q�^��7���m�����XX���+���Hڛ���S��>�����k�nV��t�@����?������a<�ؘ���~UbV���y����~��K�}x ��ۉF��?��/�}������8'�s��_���/I{k=��A0��!&^�-�U!o���?�1$%�B��gzb(��h"�VX�_��LJ�Z�����X'���t�|K���Sj�n�M�[9;�Kȩ�;���� r�e��Ai5/0ߙ�K�7�q���)+P�9�Ap:2�*���å�2qv�y�kpϜ����H>�B��n���2��H`~�e|Hҙ�S9���>�����Fx������/�+|��'�:H*�!E�ց����"��{����pKe�I� e�Q!]��! 5���hib������^���G�G��w�a�޹A�����X�h� �}�􁖟)��� X䑛��Ϡ��7��?���}�z����ߍ���mk1�N��k�kي��	iTHӒ&��'�^5H�E�.b����G�M��s:� %Q��uI�hP:�b�#�x\�=�nX)���'�;͔�t��=W�)O�#煗��Bk�a�Z�k�$��ȣ��K��� (�R�,9�-���zđ��E݄����?�#{������[�|b=2���m\J��P)?<0"/��e�CRY���Ä=�����w>e�\p�� ItgQn��յ��W=q?0�dD�d�A�AB�c�4kt�@�q�#^��noO7]-��r�<�����"/>��T��/�ec�ӾX*�,�r�������_�d�_�v|ZB��fGzvs���=�iL���)��{$���*�n�997ڪ�΃�Z��5����+J��У�%���M��O���o�ʟ�ο�����%ma��?'���_r�Z�,*6�Zc��������; ���=�>&�M?	�2��b	���zY�(��~�3]h�o�j�+?������w}󥮗Yoʮ�J���c�)b)����ו����M\M�={0��z�|:S�5|A�8z��7!�dx��ւ�6?�.CMVn�����L� 0 />=�.SU�����3'��E<���䌦O+�r�7w�@���G#1��d4�-x?$ɦPB�_5-�>|�Է�*`+���F#a��QM��Ʈ^����i"CQ9w(*��`�m9/�x����b�&&��^�1w�%7�sc��gF�ZU�]Ұ�n9rD�s�;1�Mu��٩3Э�M�To�EQ�e���{�(Y�I�ɚe�zJ_��J繁tȦ2���Z���k�J������~�A�zYq�<�y~Ʊ��F���96�-�q��_��\��}}��ƫg��g����hl�������a����\�B�*c�y�tw����Wd�*�DU�`�� �r���n��o�'��ay���/n�	m�Pƹ�-�Q��W�j�ug�q9y���8|Tn��
Y��!3���H<��)p�=="����;oK&s>/��d��[�W�S�ݨ�0*�}���}K>$���F9_��.fΜN)�!P��w�7����?Zݍ��veF�¤`���ܙtm�I����2�
g��j�������k��S��0�}EãAkMƽ.H��V���>	(A^4&,mMY-tx��1H��������B-J�-��(�fL��6�q �$���i��`��a(��c�m��ޱeJ��h�nXx0��8�0����*i����K�e`L�Р�;s˛��}��J�������-Ҍ�A��A�sBGլ;s�,{��,�tk�]s�U��(3ǀ �C��n�4�o���>X,�U1e�4���$x�xd�C?Ȝ�6ؾ�k�#�X2���xvv�Xaq�TJk��b0�@�^JN��+�Ň�^���s�1�б���/��]��a�Y�v�����/0L�o�V�5{��+ ��Q5�B��G�q��{���Jqf��'p�[G��?x�ʰyw�9	m�w��.x�.��722�yZh7�H�rBF�v!r�]|�?�@ۈzCf ��G%D�ƪ��
1d���200�����������(��/��y\��gS�7��oa*��~h��
���msa��Y/ـ)�o����k���Mµ!�@��$ꚪ���<Rsh=Y!�mm N+t�U���KջQb�Gفq�p����{���t��5P�g�#+1�=E�G33���5��x$��|�Dun��i��+P������X�/�$��S6���Ͳ��(g�8��"$ F��DU*���-Hq����?�/�"$`�{}( �q�+�A��ݾl�ɧMϩg����s)�
��1ߤ�K
�vQ3�uª�d4�aJ�EȮW�ZJ��f�������յ�7�)�H��Iv�� `>EPXև�����]�>Ȳ��y&S���=���3vD���B>�s���g�nX^'��s�p�!������G;j��#����L�EN[���L�#�2��kAZ��(�ͼ3K-O�{,�
�o�Ƶd�z;���ܸK�5k�W��U��2��<�����/�>ƙ5�X�/���ъ�P�H7���#��W�U�;����@�>̨�5�9"/>�w�9�7���He�xc�X(�A/�W��U F
F,��R�n\����(�?{�R�������2��,��aS�L���q�-K.N�K�sL��3QB��4��ﬖ��I�+
���)\�6W_,�s(�7���C��9:$+��\rv�S�e ^�	�6C����V����a-�A��G���f�?B1�W{lL�nޅ�S$>����͒ń��|��b���l�N8�7E�F�dr`Dj��dhp\��	&�jX���"U��R6�8�1P���; C� _C_<i���q+�_p�?2!�G*� �wQ�]Ɠ�`Io���M�e[�Px��v��߶1���
����}@���0K �G=j�`���,�@�]�{}rU���m��]���=����5�+�]#u��x5CRj��W�z�$����m��7(&����=��8,��?��99za�F�0�$���4+���):�f`q�-׺M5p	5�kd��" ��Z�Y�IT,0p��Ldy$�pZ�����b���~�2i�\U�.��m;^%Kw~B�@��
��l#�����Չ�6i����z�^� M�6#��(�)y�sCX7<�)i�xK�(�o�,m[�n��s�7 ��O����?&#�gd�e�a�vݩ��uɖ�$�}���F�{���ɓ�(9�A�n��\�Pi���ɸ]ħn��|��A9�o@Z���Cr��QY뵘�]W�eg�v��Y�������b!2.(JM&γq����ft\|�Q9q�Saz������0�S��b�WK�D~��7 /�B̦��sݱwp�3��Z]��7�X�Xj�E��T�rH��&��3 +`�{Ē�i"B������%���j�=ts���jM���������g+d�c{΁W�q�dEn3�O?;�'��5�6�
�p�Qw�]ڠؤ�"��P�7�U@5>H��,๲�/�ܾ�f�5�[C=�QsT��N	�0��QHW�~Y�z�t�\���!}��gJ*�{�,��
?�O����
i�����^�1F�v���E��9t� bDF��c9�p�U�ăX���@�� �M-kaIe�HZ�+`Bpۨ��D�	�Fq(5���+Fw٧���x�wP^qǣ1u�RY��ԨL�k�*h
P�!��(;��&h4�7,�������Qݰ�*�#LM 9Q��B֫P�Bp�V��{�~���8*��8t���&P���[�;n1�^7���W��8���%�[?���m��u 2LL�9���\#��5Y� �>�\�����
�	��ƂR��q\�Qms�S�r)�{��4��:�&�U7U�Z{��T�3U�o�^��R�0��]����q�Q�a�(&-^�zJN�|H��B�b���Nd�U�m_q�Q�"�И
�Оֆ	���wD�{�}A�B�l*O0!ߔ{�6߅���0�� qD_Q��2��腡���b&�>h.c�1���i -M��KS;�$�|���}����2��|S��B�T�]��ь:[ 2�7������	<�V"�s�a~{Ж��^�ﻀ:3���xs�[�D9,/����/�Ї��k�@|���<�F�ЀQ��%ku�1�־�-���s�;a�a�"��^���>ٳ�y��t�x�n��޻dͺU��
�ڋT5렻a����XS9�	���\]w�\�)�ٻ��'/���t���f��
xŔ����..�#$�I�U��10"c8���$�&�4UV1\�#��n���.V� �Ts�]l�ht-�ֹ���x��`H��2�JU	�ҵٚ�u��c��r{ �b���\��l��Ti����b��W�l����nht��RE�:*�p��5��`C
���i+�q��f=���Ъ=0Ks����Ϣ �	�����E�R��L�tipn��8�	'
]p�i�=����B+r���9���Lhɇ�8 ��T0 �q�����nR��	ॵ��PŸ1��p�E�SF����	�J�E�~���3GrǏ��keӆ��G��'�z��c)
�"m**]O)30�Y��_� �vy��7�U�
��+�H*�X3�׭��|�A�q�~S��F�	T���Ȏm륹1�A�+W.�eK���2��nr+6�G��e��Un-O��*�yƪi�هQĮ�8+���Ĺ��R�b�M�aρ���y�q:Pt�˅� H����(nhM��ܤ��X'�@��M�/Z���r�(��r�M�;e��,޺�g\�W�2?e���|�+h�6<G��Z-�SD� �,I�eJ�t���x"5���+�l���Xh�,b(�8ɀ#	�f�o@�M�%#+@�D�����8TKc�uM�͚��X4��Sx����^J`Q�qG��pcB7�����M(����^�8��"�7g��]�o�p8(˗��-7�(k�vHcc�Y�$<�;~��{�YN�>¾�T��l��ڻƐ�._�D>������/��*!	iEx\.\�(o��O7-�<�p��e7���x.����M�R�9��5�����	L/}^JXhL �r�v������Y>Y����\�1}����6�g�e�G��ݜcֲ���r�kSI�wU����Z����J|Ȥ]�X���Z<���!U�M�E<��<"�hz�TV1O̏�l��8d_V� ��1��������29�1��J��(�f���i��[N��!���Tm�e%B�¸ .V[�Ќl�4 (�c�O�Vd}Ƙ�#&ZRl.�2;(@J��;��k"���81]��-�X������ٝ�{���9��,A��)�un~��:�+p*���A�L1���XؖZ��� >�.L�]��4Ț˿g��Y��Us7�x���R��l����X,��*��L�'~�P�=b
�R��|JKo����I������8����'�~���=p���tXG6�H�O'X�\���j.���7-��0X=���v�c}��6��uj�[�ʶ��i��(����H�g��.���
��	R���`�c�g�p�5`wkG�|�~P� �{`$&?x�tG5�_-�Y���G���jFnYKW����0$���'��A�f�87�?+��e��Ϊ+{7���0�l3�ɧs�#� 4�������X~� �Dq��*��BA�ƺC�mJ�zՔh������E�%涅�J��[�S݈~�~̨����j㫇9���.�M-��&�I��63�}Ph��bǔZI��bN�#Uw��ޯ�����xLR�O�4f	E�Y2���Y��j,TZ�s�g1�m�֙�c���������>�u��� ��ڰRB��;�J��YS�D�
9z�È����ТU,�ĸ��B-c�i����[W;����1y��n�h��ݟD�UC���L@��A!Qk*>X��'�aC�H�V�����pnw�m�X��0�{�ʯ��<�	�WQ��-5��#�J<�=��3���B�k`5ٵ6$M�H��3�ܾ�Iy�tT�HEmUK{C��]jb����բ�ˋ"r�`��M냲f	by�myq�(�M�M-2b�S�!õ@٩ydܬ||�z�l]�xPāR��#�񩷆�>�(ob��̳fB$e0���Ta� GP���g�]��RC�T��d��S\B�d˵6�{�sK�����DlX~�?|IBmK��C	t�B� �/�jg�*�+]^f���(S�?�H"�΃����H��<�?���Wk���vqF@4�`ʰ0il46L��X
}nw*c(P��I՟u���֬4�s^�
<=���p;������ ��4��B��Gm�v�-�2S���w0�������r^�{U!���q��H�Ԋ���n������:��55��`����.�gFw�V)hI��#.M���X#��3vF�6�(GlZ��E�����yFѠ|����3S�V�Bĭ.��i�l�u�Jy�ٹ*$HP�mk�؜��z!�B� n�t��戵�g���H���Rm��3o���x�AK�L�N�J&!`�Tc�1!p�ur�F	�n�~�W�$���}�Rٸ"(� �v�/.��B�<6v �����,Q`���%�<j0zUI!y�=�d�
0棛)
����٩�2=6!mm ��<xS#�`7��ڙ�s�_9��7ܲB��Z�뎀lu򎎟�DoD-`�u>y���y�N�y��9�m�wݺR��hA�0R�_�>%qЕh��9�	 ���Oƅ>x�rY�fuzc�w�o�����@Y�� \���Ƌ syKPv߰�A�!��ǥ�+!�7�,N6��q5rԀ�jܯ\�8�� .l�8!	��7o��h.wR���0/Y�(
�k�7c?-�`{0-��΍��-�+tQ�`·�����	H_s�#��b~�30DM�d��r�&�
qL�8� iɰE�ƪ`N6�+����j[�tהk�c�^j��/�)�湥�~�g��eL��ThrV7���X��� 6�G�?�l#ߍ�b_s�������c�Q��q f���u�������H ���m�7s|� �z���bFw#�疙�V�%g$��,Id,J&-^ǅ�۲XZ�'S_���^-u�n�Rs�z�ހfX]��d�%8� �$�3!-M�҈"�M� ȬD]H�x�߽`��,&���:8h �нV9u��_+B�r�����ҡ�oX�c_����"�|*�Ǖ�5�E܋�R�&~�8�|ǳ�Ha'��5�A��x��и<�'�<c�9��J�nx�.��� +�ߺ`iJyv�E��3g�sb.,�lٶEn��1X�f ����H��:iY҆$�Uxe�>����>]_L�_�j�lYO>,�=���jp��S!#3Q	5�I��ټ���I�� ���R��TT~��e�2ԕ��s���!0\Gh-�+@��2�����]�9�H
05�,�9����E>d��rV?��H���⇨Z
��Y�`���R_ߐ1�+ۃ�ae���݋ L���Y�l/3�þ��h�]��:8���=&G_���]wHW�.�pR�TUN6��$� [�A��cm������ߒ���rハK�������Kq>���A$�T�E�r��s�-ٍ�AN8@�:�Mx$�4�0��|/¾"3>KP������X��m\�d�&m��ˮ�L�8̯���������k��Q��Ij�@��n' (l�t���6��ȋߜPC#c���>��������>l�g� yZDV
��nj3t1�� ץ�����Zz`�c���AN*\ ��"n���Y���;;�C�F�^�4� ����J�e��Qˤ`��M*������U���jb�'n��,��r�d5��=%�4Vk�]��y��0޴� :��m�1y^���^���ἐ�~A"���ͪ�U�aC�3�wV ��iqH0��P�T���nW�5s��
�Џɹ�^���n|֖��1�1��d��!K��.���r�\R֗�h|c�#c����s,��;�����p�g���Ӳ~��(u�)Ǐ���1�j�'������1$�5��O}2]dX���u��� ,!�.��Uy�8�Ge����,�j� taM�&``1]	�n�E:	��+^C�i�`2i��\�M�t��k�ֹI���s�ٻ��1@�]�}����9�4���o>�'���il�`�f��L��X��d	�ܐy=�e����=ؕ||�!� ���np_��b�6���g߁�$4��[$�0_�ύ�R�D��ÒKup5n^S���}k�<�ԓr��E���Xw��P�$�,/m��\-=�����ml��?���B������<�l+*0���r=�C�5�u~(� �|���9_�RۼFF�H�"�H�]2z�+r��!ܠV�v��I�q1�h<��<`�k>PdM��*��ꬫ��*��5s��4w�Jh(qh�`y�r��Y�#U�G|�vY:Q�}ps��_b�;��[O��͝`�߲S��;^�%,���Q�t�H�b��s��<��^�$[7��}�u���ȹsg��V%������C����C+4�N1��~���	v��Wn]�B��'�z���}�|K���h"�R�Z���2H��qV�/4�ܪ�����%��*{�R�ŭ���O7�a�3��9eY�4��z_~_�s��>�%�Dfv]-iL����.�k�Q�J`H �}P�>tzX~��L���%VLC�=�c�lt� 2����򣳰~�� �S��p�\xI&�O�����°�n@��_��/J��O���j�9��_�5 "m�,,��{���9��R���u���&˽E�Ȃ	�jy�'����S�y�G�1R�C2>�2'�>�.��h��~S���X'�&����`�󹾘�j���� �H�}�3qB�����dи�L�`�:HM��ϘR��o�t,%�qV�9�⼋�\�w�Z�������]Z.���̞�>���x$!k���#kW4��eʚ��wrX�8�#!(P)���K�X��>�������կ��9|}>	KUH�Nn�i�r91>�Zĳ�� (#���[_����[�Ɩ"�	�# ���ʞ0�݆aٽ�W~�w����N�:]+;>��X;��ߩ��nh�����o��#���w��K�]�qSHs.��N�2��W%�]>_��d`�.�^�\/)�ʴ��~:R�edY�l@�-ʝ�e�Sf��V�%�߳�7sϒ��T�p2�+����r�bKGHn݌�Π�04����BN�����Z�	bul�g�3r�Y�U��R�'s��h*vA�:O���Vy��3��]�06����ʌ����db\�䵠}�~tIvGr�'��6{�:���TLٴ[ ���G��6S�+Fs��f5�5"c�s���'�����.'�m�q�H$w��Xlt�,4@��t��#�@����@���c��8�� �
R��;����2�Aˑ�֨��C-%>��jL�W��ʻ�F�����ƭ�9C��gr���YU�)��9����3ݼ�Jqd�2�d/J��č�AS���9�*ܙ#�܊����~d�9vVZ�p+�L`�C|��6���TQD���AUf��tDg�Av�ge���˸�K�[�|b�D��c@����R�<4�2,�n�> %�O	�*��K��1c	ܩL���;Sp+P�c�����������{�6S
.G*  ��Ӈ h���}�D�����T� GS�P���� �s�L��k5�5���D��ŵ9����c���!Ȳ�#�D�%�����Ć���o�۹H}�w-�T�~H�����b��+�����"�뵩YV��e42)_��t��I��IpZ�Ԡχ"U����7��w`���Q�6n^.U�+`�4�r�$�>/�_���wI(��dtd@]�}�S+}3�q����5pA�Cr���I(X�=�#���,]W%���+Ɯ�$�{nZV!���r��y�� ���^�Z��y!wK}���>&Χ���108��|r�Ai�X��r�pr��j6�&[�罷'�m1׋Ιٙ����l�b��L�����Lq,��m�m�EY��<�����S �bp$�p��!r�@�7���o�Ze l,�kcn�1d�e[st��$ۚD�����ac�eߋBO�b���7��%��*��	�*Ux
u7�.:�%�M��8�۸
B����G�ag�E9s���ZO�`t�� *��"D�F/^���L��HE��!�(C����y���ym�N�����,Y��O�u�M�m�*�����APx����|�������h�7sɾ?�9Ғ�-�a$��0&�ǁ�By�"��Jz�
[�`����(�1{b��~YrՈi�bC�b�p#��5�Tj��^��=�H:k�9���ՍF"D��ī<���D��*����Q	���dA`���&���M�7�ǚ������9=&�Ȫ���Dv�0-d �xݓ��w/�(#�* V�H�h����Ͼ�/�:��?�C��L�
����Cg�囯1H��i�3r�E�TA �����换���0Bz�����Jw�Oʟ?ua�C��m�:c
�t���WQ��4٣ ��]�Cx�R������s���>�c� �q��P���Xi�%E2�����N/�;��Aiz�%��Ij�l��q�L���o�7e��[������y����GAl�x��GPY ������{眜~�K��A�|a֢>�c�j'VLE�̱�ճ��D���)+&�$�ќw�^�
��u�K�V̢S^�f�=K���t�}��Ks�~��`������ZM�ٯ�,#� DG�]�5 S�b�.�p�h;����xZ��2¨�>�[�ٙ����b�* �Cޔq
��SR�1��>�;Y��ԠhGbUA���m�������-4qT��w��P�@g���� A}�=RW3,[֘s�|�����W�J���ˑ��w��;	��:��_���|����wބ*�n����j�Ҏ7�G�*3� �Ljy��M��5��:Z�W�|Q�+S��s�m�᝱,L�(�Y|�o}ݝh\؅���|b��֎^�ݩ��ڇ�Ԍ��]�-��<Bk#��������X����dXsٮZ&�n8�zV�wv��ה'����jyp�_ڑ��̻����ݰ�e�(M{���C
��\1�x�!��m6��hr+(�f���i���CU{��}iK0�Ě�|�g��U�C�*Q�fcm6�=��F���Qc�Vk�q1�u6#o���Nb�[���UA�yH�ʷ^�����&�xI�|Aư�\�{��B�t���V�5�\쓣�.��z�� �kP�e(�\���Z	����_����{�2a��`Y��LǾ���b�k?C �8f �F*�ŷ�����1��w&�c�$�49��昩_-mKNI�Oˊ�l�Q��E�}0>�/V/Mko�5�NAލK��^�_q�e�6q#�ܜS��܋�2z��:�� &�]��)����u�,s����`��C�Q/MFe��E9z�< �_���~���#�lc��Sd�Ӓʙ�R�cAJj^t���
�413��L\
��et�����;c��[��K�/�z�ӭ����`�Z.2�h�i���Z,se�
���|2R:��A�Nz
�jl(���������p�A`�8΍��lk��u� �n�38� ��Hw@K��|GW}{=�Ĺ� � k2+�8�Q���K�ĔT�y]
�[K�Xp��� ��H�x0�tgi,u�|LƲd���1K����n�z��m�gӥ��xn֌�����~l��_j�����_�/��X�Rٯ�� @��:v'B)�_pFA���!,��&�i�@�d4����)$�xR�Z���k��-~�{[�b���l1�B�1W�|��qY5	�U���ڮ,6�c�J$�=����la�%�/�2x���T�,�0���"���G�g*�/16�Yw�Ս�&�϶�d{�>gf � ��>�Kս��3�(�ΊH
"O@Lᷥ%�f�ᦟ��m��,��ڥ�E�Y�sI���~�'���l��ؠԷ-����yX~�.^q%z`> �=�e��%T��e��M��!$�S��=Q�d�[��[�o���@��F�����S�6Q����i���Xk�7���*�N!	 F��.$�	�94��
Z�3��٦Xc���������)�ݚLYMr���0/��h��/��f��@��4g�4IHS�
w���S����޼~�����?���:\(,�8G����ԩ������ޏ9��֡��t�9�l��o�%�fH �6
1�S���tB�~�G2�e��ݻW�������?*���ú�g<�2���².,t3|hf�ۄů�9�$�%����h����&�ئ���y��c�� ������ ����A��,_��5����Z��<�k�-f{�w�A�͍\,k�d���3����`� �Ϊf|[ �`���*�����[���>�P���s[T�=(��\r*���5�o
e�jo�.f-�*��\�DW)�ŷ��*���\/OU�K�.^;�=0����Y��^\t2m95�K�X�ȹ��ex֟*��P���Wߔ]�>��v�ʋ�M�:m5���RAH�^uJ0j�]:�'��qq��~�L�������;���bs]�
Y|��|��ԍ�Yx�� �vd�>�B��Su����{�ų�=0;<�J�g�Z	n���3Й�A��K���$,�s��oη�E���`ɬ���i���7��'�/���Ê:.��o4�b���?����lPX�4.�5���k��g#���&�3�Ӎ�\s$�e�*�A�Ȁ��A�����g ;AA����5��[Ғۊ�á\(o��8�]�6�����t�y�z�Ip��ٔ0�j�p,����(���vб�8��������S�9�k5�w�,�hh$J �g������af/����F]<�����G�][=��:Ι\lӰ5fh��j����rc�Vj�t���݃�����4H�|)ب	�uO��*�)[������x�(��)�P~�iEk�Z��Yƍ�ڳ�1J��B �9;/��|m�㲱���{@�2�Ϝ'�S�m���[���Y�p�c��ufM�QM�Tl�V"���1{Ιl��ɼ�^�_��~�����k,S��]��~+Qf����~.�+-�~<��7J
k��-��a����:��La��Uo�8��H6�'���.���5	�>J�������xA~΃�i,�,* �?��Vό3��cH�H�o�'Ӆ���~t���nSZ�L2�\%Y��b��y�#,�1e�@#��,����� @꿕0�l��N:.&�R��#\�A�&��Y�\�h�k�p�-4`2L�$�s,���C̸���x�#r|�{r�l���d�M7�/$���Vj�v������Cp��R��pCj�����`+zP���)
-��l*����w�Υ�l���C��;E����Q��I+5e�*p�!i�9h�7����v!���͒T���ƍuku�=�j�]��"��˅i� �J$�m�cn����`	�V���.;��f�/�^ރ���&f��.��|���D�44�ȅ�J�K1�vj�nD����p#'ǘ=G-g������ޠ�p�+������L+������f�s�� ���iB��d󮙌?�(�Ni��iY���魲��N:/v�g��Jp�OK��Mc����z<s :�dB.5��$�Zf\�kp��V�:dP*f��xˌeD,)]������
9�9_�K�T�s��FN�^�&n��� �y�X��Ls�I�Y����c̞��}�T 5�X)[�q	���Z��6���~[A�Y}���X#�j�/$Ԭm���6�}��sߴ���SHDY��*���f�)�q4ď�a��CNs�2}��`n#��]�6�_�V6bKs_^7��;�־����p%�yO
6�#�7G>�����>
H-�L��+&vj��.��w��f���J�>C�&5.��Tmg��0g�B���a��]���%�,RJ�Fh�r:F�A�� �T@��NJ��:���X�:�;S�VN�q~c.��ufO�����V�fd��m!1�Xz��Tt���R�T�7�ߴ��~����<�=gg��&���#r�!�Q3pY�XҨ �T6���
~릐�ioE2�^y����k�<)�]�T��?/��y���������J>M�**T�.��Y`i���\��,�WT�H���E�e�֏��j&ƣj�%����|0��Xҙ���a5D�d^�F3/�pm5�4��P�ŦRn��"�P/�w�`JϤ��՜6��Z*�VC����9�m��-7!�4iWm�e[��	{����mjW��
���\�wP�I�� ���:J�X�p�$ۧ�:�ci����o-����Zinn�o�
 �y�ihX�*��pm6Xl^��	�������L���Ta_��&+�j����c6(�B��5���e���	�lw[���q�[a��V)�O�8%p�`/{:]��O��VX��A�4�x0���c�Nv�Wfe#Pn�d�����I���J�J�� z��@���@�q,:��vi�7�+]���p�ƔZ�U Ƹ{͡����f��Vp�2���6���/�g� ���G*-x>�=�'�<f�'84V$���D�}��&ZR��$�$@C�$�3^ՅF%>���3����������t_�T"�If�Yr�43W��{1
 �w5��7O���oW����e� 
'V�'(#�gP^?4$]C���je����/>�Yݛ�f��{��������	�@>3���F���O?�^��kU���A.����	y�8y��2J������S�wa?
ǥ�u�$�����>-��֞��u9K����/w�`��6;��sǲ�bxhχs�2��Z�=�)���d�:���V@����H� �Rr�uC�uF�ü;��GAD�h��Ѹ��om� ��Z�o����8a�h��X�|)45�*���"={�� �3Ys�
�`K�#E��]X�%{#� �m���'�%�l��l��֨�c�S�:� ���[�2O+~OE��
����U���������g��5`;��Lц	^)~X6��f�e�t+Vq/Γdt�8�����A�Q���e��Q��q�>��2���`��D,M��7�_���6�5�8�
D�a�Ba�u�D����ͩ� 8�Yʷ�R�Oˎ+��h�cj��e�ʙ&��?9��f�&����vǺ�9�In5��c�H<&O=��pe��܆0J��K �	|���S��]ji�h?�9�m5���o���7��7u7��7�2�O)v;���d"�}�Y�6$�-xXxE�Mp�b�oc��/���>ؾrR~��Wd��y����%� ŗ�V\f+8E4�W�/S,Ի��Ο����Lg*�	'��s��8	�R�ys�%n�y&�n%���ǘ�3H��gQ�b�Kk��U����[dw -c����@7.JA��-\b���_�=9����`)@�M*7�hB,��$�>�
aS��lv�U�B\�:�,8n�ӗY���0b���q�3�
��D�Na\�ʹ��u�ǆ3n�>`{�{eKP>���O�Z�����dwW����Y��cpn@�!�4�8�x��9�D���'������s���ɍ[:d��ذ1�-u߀�IPh� �$`�!AK{dǐ�A�ej�����:|E`�i����j�&��)�p��Zqp��\S�{��և䐍��˹^ %N��~6e8�X�ż���f����X9L̑ӊ�S���E�[��t;'�g�U���
�sYKNk1�I7�]s5��c ��UHgl����_�����_7�y�����o�v���3��U��7��j�n1�ԲV�5��m�n�1�k��K�5j*HEۣ���C[�թ��>���(����!yso�\��)C�_�5���[�A�pƛ�M�Y7�{B��mW�x�ڶ5`7��ǵ���
�5�鮘�6JkP"�j��ٸa�0��`�`1�|<;���bF�f�Xs�h~j�w�j$�%�q%��tOR� P����`�9;��F ��A�9� �`�Cس����t�v�������P��RRe���U��QLk�~L�`T:ƭ��&n�9Uh�>�r5�2�c�[������M����٦=z/��(���;ҽ`6AV@�Y�	vk�q�jX�3�p���:e��LV��9z\��%1<<GH6�c��<� ΐjzU�������<ǡ��/��H���)$B$�8V��vEP�y�-y�/�u�5kW�ͻ�ɪ����>}`�} 7�Xctm��$O���+�7�V��` "���l���޼?�J��ay�n�?�8xm,Jģ���sF�B��P@!�����i�F)4H:�1Wx_u}���|o�J-ꬠ-�]��`]��ީ�f�Ŕg�H���F�Re=��D@����
m~&�t���w����3��q���%9���P�J�:Q���ȓFpG��@p���ð��)�;���вR9}b��<�6��1�6�[ƌ��Q��R�L?f3���BZi��X�Yv���433��F���&����@N=�}w�x�l�夬Y��r	+K��wm��?�����K+����Ń��-Gf_�d�4n> SA����剗Ql���.�Xx͍�#��1O(0m��k�����Z��{58��c���?�Y��6-���2�M��ǫ�\��	�!� I�@x�;�Z���&.'����B@�- �V>�U�>��l�hY��S`Qpf��T��W'I�Q��d.t��
� ��y�}��D��{OZ�~]J0�)|�֢��(�i ���n~g�wmm@�6w�_�)�q�����ȑC�ՅRhk46&+�!�VA�y��@ܰ~�싌�t5\�q�b��f�>\ѱTv��"�>Μ=�R\��tvvJ��yĵaU�JKs�t��o�"a���>}`�G�Y��h��>Ԣ �]��:|f�75]۴:GZ���y���b��Q#mX�������I�V�`8y27�����k�]Mdȇv�-'�ؠ)�y�+8��j Y���R-E��&e'x����gk<���t�qcg�Ɍ^�{*X��X4�����F�[�P��%�zVJ|�L+2s��t��:����_���x9��S?x6�RE������W�/$ê�F��8!���"�WT�%4�0�6 �o"��U7JC]JȰ�[�QY�Cl��А|s��Zۍ�	"c�VUP�=cJ�-m��JC
2 �����c�(�N�a�P�˥����M"{xY�_ο�
�tvj�ើq9�ڷe�Cw��p�r����I���u}u5�`;�43�Ԓ}�| &ޫ�z��'[�5I���Bky��oCy��@�M�<8������VV'��ވ��Z����J���u�<G1���e*<2G��(�(��nd�5)�V��ka���9s=������T܃�(��]¢���
��������~�y�����>XD<�yT+��x���ˇ�[���u��5��x!\K�7��_��_Њ����=I��Xd����?wQ�~�D�ǱA1SYSPFr����?3�v}���V�i��n���?�|	Ndz~AFn,BZ����7���_d��Ur��Q0T��m�{_��U��J �r&�d�V7[����s���N�g6��!&x!+`D�TS����BY.�%�Tkf��5;@�^#l���2��q���i紺�^�C\Lx�F��ɗ���Jy�T���H������?%��(��%HY���O���"��f��(\x�ޞN��?���|�N��]9����{�I�f����1�<�&*���rཽ
�W�D���ci"�ļ׺�hw�	s�.g�!F�P�T:�\.�ĥ�['��KB+��č9.!fc+����f\�r\/\��H�� L*�%��.FМR��A��Ğ�-�]\,86˗ ��u�#���T�(�x��<��t��#��<*����8�7�-�cg�Q?���|����c�a@v�jQ������@�
��ٰ�]խ���ΧXa|�?gf3/��k�&���u�I1Ͻ���ZBep��iiA�~�k���hœ�t)�y�J���r�d�
��n�&�b�ݣG���X�,e���!VW�#i�p�87��Jg1\g>k|�a�V9���r����`�ʶ����*#Y�K��|kJ�֤s�H�\�
�>���3�Q*S�%BtQ�UZ��Di�<}H�R]��[�O�xD�#�mI\}n�69���~ܘY��0}J~�Mx��ڇ�%�7J} �6��G�zС*�h�U+���8�8M͠q������r����;�8ҥ_#[�l��{(��o��y�$� ��y�������pXV�^-��Ѳegީd��=x��D�X�Q�탭�r0P_�['���2����QF�Ț&"�8ZƒR�t�T:��� }������I��вi����Wg����2�D�}�o�V��v���'eG��"�v�NVld����j�duMw\z������]�	�����4���&�W���ن|��^��?
H�rz��e3i��o�����t"A��!A�`Џ���$]<�ԘŒ �Kq'�<��Z,4~����+���`�UƫP�O�솪����(�l YK��ʜ͌[�W�C-�\��8&�d���������;vۮ�%@jw�!v�AL�5��@�����?Rth#�NP��Zv�E0R:������1 �|f��X0\%�e� >�A,ޫ?��N�.j#��ѿp]�wR�D�rd,$=	�,��l�Ph�k,�֖�f�ƺi�N��<�n~�-ޗ=�bĶ����cO���蔌��Q>� ^E�`"A�iA²f,Lt��Nii
����¬�ad\��4-���ukr�!2����P<"up�9Z�B@��� �@�����2-r�m��a{����"�G�$жS�Zd7^6`�ܚ���C���((V.k��7���:X��<$ǝœ�v�Nϖ�����\�W�\���_�͗�i^کZ�E�O	a�|�w���~Z�J�Bg�F��ʘ�1�l�R :�]v��=�)��Rm�L��h7��Nݴ��̦`z�����9z-7Kŵ���~5��0��U12�y�DΛ8�� �	�9�n(i���\σyo��}C*2t�)x"�#,Q��1.]�Y/Pj-����~L����y84�؛�e�r����O �	���W�E���9�b���p��`-��/�{N-O�d���:
*��)s&@VɄ���q�V;Wo�ٵ E~\ҽn%t�/X)KC+�L�]��>�|m8���-�|T��J����fm�,6g���ϸ��8"KbRۺ����a�@��b
)�z�2��~+,��'����>9<�V0�1U��c �o������ѝY��Dk[��NXx��O4��m����e�?~J���G��༘ 7^4����s�$]ouu����_ze/�����s9�/��x�G�ʷ�ɍ12�ѐ��Z�JZڟcĥ7�(�v���c��A�`0��u��d�g�[��|I�m�yݟ9�i�;ɀ�RB�LOu	���?U�q��9�3�l��ֶԘ�2����ĹݣIB
B(�MqP�zr�J�J�
v�� R7}[�Ϯ�׶�)�v7���f71 �N���t�d�!6^ܰ4,�� T�ì�����f�R�_Ǻ&�k�~��s�Yȴ��f���t�O���e[ͦi ��@7ja)U� �]�_�W�<d�~`�=cQ4��� ��R��o�b�#i��A���ռ���u?��R�ך���]�v��*�m��˧`�A��&� ��%�X�5%������ K� ,1�.5�A:�L��*�����<%�J	i]�F6ߴE�A�?x�^��01Fƚ6#7�f^Ը�2_�s����[٥�֚l���S?Θ�	����oe8��I}k��pǮw�+�fV�s�
֙���½4�r�i>K3M��Y���iт⑁�Qy�=&�8瘖U7�Hpi�!���'�}�p��9x�7����ޓȣV�!�?)!_ o���+tp$"��?�� �gѓtuɭ�I���(%��m1|Ι��`��_ϖgn��y��>�h���;sN�K�Zn;��W0�(s��$�'�!�<Z\e��*�V�f���0ɰKВeM�;'(*m�!Ӡ)5h�|u%�y��A]���[���L��,�S��(�{{qZ,<k�op�2g0q�[�����7�etl\�;��9
Ic�!�|�ȰD��Moh�*��5R͹o`YMpG@��}��e�y�1� �����1��u�(��<���kI)��b#�cŮ�`��̩l6pAH�!dXnO;>c�jƳn`u<c�����k�T��*پMқ5^��p�T{�aU'd��[e���=�)_C������-�$�TBSg)�Μ�G����0^��Z���z����CǙn2�cݱ��QjY�� 	fiŲ��Nx�������[���p?��F�S�Y�	�-��.	0���nbU��2!d�����T�Jy�j�7B�
 �*�c�S͒,~��i��`��C �M�P�8�	I%gxx����n��0�h��SFY"��wNTO�L�So���p|�}�n�j~8���l�u�54!?|oT��k0&p�-�2���Ӱ.rne��y&�iZ�<4"�󇐸�F_�1L\f�̯Bʔ�uA/4���?yF��+e��M���|�Y9�/{��TaI����Ӭ�����`*�2��̪���,�U�e;T�s�{8$
iM#���2��Ų�U�D���
Ztˊ��)�f��'���8�'i#[���b�w�U2f��	ʍ s�~j�hod���<� XP>J�l�t&�5V��n�nQ�.�X0L�X�#���rۥou�h�t��dx�\M=�	����z�''߮Bzy�lܰF3���@vY�_V��q�Q�����ً
dR�3f�������!������]yj $�ӭ�4M�����i&s�!פPuc�,9��l��1�B���#g%X�c�ϸ��A�C��|_��&��L_�������l�Kk��a��J�Gq�1��v�-´ta���(#8�D_P��!�D,i�,7u��1�J��,#�r)H��[�u;e�]���0�n`	c��{�yL�kj��T��U��p�;=*'"X�l'�H�i�f�d<Y�\�b���qYJ��N�{L�9t�Y��խjnV%�A.�G������LJ4g�ت��G���T"	D��rq 
�q��S�`��B��N%���Pf`���Fpbקsޏ�˒s���w�#�X��r�<S��y_[�7Y�o�Eyb׮h�عw��g�R�;vIݶ�q(�$��%��������j�»�L�r2��*}
���X�I���&ل� �^ۼ\�*.�XE@���`��z�n(�!����1x5�{����s\�p;(i]U��7
���B���:\6���`�󕯑^��Ԛ�$��l�h�FU;�~�j�kʤ�	��#SsW7M��J��=4�lה�4�Đ����00K
$�����R^[Pc�қ����o����7@��7
����z�L����������Gŏ���_���;wFA҂Ts44i"��#�n��<�E��|���Ո����	�W��m�bDd�G��i-�@���A�|��:*'O�լ�qp\���}��1�����4l��T#�v�r>0��`3>����>��c��.�����gu�!=���0�L��r��Rl�x��1.�Ej17ɞM+���<�<t9�6�?�VT�v��?�ғH!�}3�`>{n�	�����S��:"���_.tv�:�R�o�rm�@��2���6
3����"C���;����Y{k����"��uYxs�7���K�ӽ��O����*�MC�k͝�̤c좒�|����6hĩ���`ڍ�{C�o��N�UV�Ðvw�n���)-c;W��^�%������ߕ���?�e�L6�'�O/H�n^��zz�� L�AZ�Mm�h�vW�j����ǣ.�< 5Άʸ������i񅨉ҿ��,�ׇ�qM,���~d��ɑ(�����!�X
�'��0Ú�7WiP&6��E�֑>d8���	�rjT��!4"W�\&^���%N�����ycx���,�Q!K�kZ����k�b����w����R�IH__������=^�!^|�z�
��!�YJ<���	ڒ	�oj�GڷqL������!,�^[W��Q^	 뤺j�j�����.3A���B�
}�M[=9k�����L|W#uW�/�N��!��ʸ���ȅ��="�-��s�}��76���%�/��q���)�v���Z��w�q����RW�V���i�D��|���*�@Y��	����|ʚl9s$���Sf�������[��ץu��z���z�]�C+��Ȉ��o�����k��i}#~ꤽ�vS���k��A�ک�˞�<ɜe2�L
~����g�p�_��7*�ؿ�},�g�٨|����|�_��˿,x����9�����'uX�Tj�i�S7f����F��w+{.�k܂�� v���w����o�,���z)X<<>�->(��#%�˘���,��Pᮦ���.���0�z��.Y14��ib��h�QK�4ެD)�����:��{`W	�E��woǽ�%"X��\�A���g���S���Ֆ��(�#�l�i�4-mV����B��|p`H~���g���̱P����e�֎T���6�d{^xU�gp�L����?�RihC�#��p�b�cm���w��#r���>�@jW=oN�s-5�Ҥ��F6���*yolO���&;#ߝK�)�Q��`6�AKvw+��{Q���,�U9���]�4�3��h����d�\�'KbQ�NY�å �,/�n/�h��%�k��2���~�3�r���rn�̢;v�����h����&8&���DF�p>�����*(W�G5�����Q0\��K�� +�$�Ve��<-ybZ��_!�����1D�
�2C��9f�w�I�%Q���)i���={J�"�����]��+t�9x�h%n��5�2
�R�� ��ODy:��9� �1F��>魆��Ȅ�!|�W����v���,Y�04����Qy@"5���J�
����S�-KV/���]20N��.���ՈC���&@�1S�x�҃E����������¡+�em.��\�D� @-N��5�	b�I<�4��(�4�.</~l`�oLl�EW �����zC�P7N���SV��JV���g��)@p����������n
��s�����%�kG�����w����\@bL���:�м�K�F�b�9��{���r�0��ǌ"�-��'��;,���� ���$̄	��ęC�H�td��j^���};���w�w`L�ݾu�����aG	��A�|�~RZ��$To,+��n�:T.x��%�nM��L˩h�LV�I]C8����ZnjBj;�f{p���WW��U̪��932Խ_�'�];Z�B�,�,wc�e�;Q�m��˝��ޭ�� �93��ptE8�Z~p��2������o�R�8�}���-��x ��%�so�E���w6�Ⱦ�x
�Ny@�����{T`�4n��,k����ɲ?(��U2 ΥB`��H�3��aD�W�=�������>&�N\��p�M�%3��Pܖ����⹅z`�+��>�F_ee�Q�o�����F�� �Y!��5�B�6�1̻$�i&}��g�B�p����
�kŲv�Q 2�8��T����N�K�Г-T��rڙRd5ƫ��T��6Z��g)����6��0����}��Y<�2� eM6�i 	���R��Y]T��$w�";qo7<���+�Z��w< ���Ru��*�y��,�XS+7��l�z�ύ��K+��(��Hp����*U�B$���/�o-F<�������(ua��[��/.��#�aYP�B�ƹX�her�W)k��!�5�����\�\�JD�u{4���&�4���m�뼗Ql�A^���
�5�!Ӑ�e�� o�#H1t�N����a�F�%`�fˊ��ws{L~��#��9IT���G�$�Ym�����Z} &G_�;�x�Gӷ}7�ӦOK$�}��\�9L�|�| �������%چ��sF���G���m^"k�U�nڡ�
���|����ìW��F����&�9aX,�]��v�wH7��<��s�=;�,�@�?�Fc1�m���ܸ&�\L� ��������R`� �:z�8�Y����DM�����6pZ��ie���i�-?f���HYdx��Wٸ�QX �W���� \j��q]�!ܼ�}Ҷn]�/K$ǘn�>i����K�[#��e���Q��.�"��\�����A�ԃ��f���em��t��Jq֩�
p'&���D��Q Ɨ�rcUg]�$������R�N���DY����kW0���ƌ��9���;��
��#�dX9�lK�ᗲ�Q��Z���&dc���KQH�^�=��
L���? ��3&	^^�����z_���|E�����/��Q����7�k�����v~w��x�lz`> S���r�ΝG_C�����3]����V�l{���OW����ScL�������rL�ZB�V:�5p5%Bg�e��5���yv��v�y��6�i�~R��E��5`g���ש^��E�&�5��4�{5���D�3�?�$�,8t%K��v	MO�9����y����2t���T������f,�c�4f	�N6X*�@҅ ��8��WYH�2����Y��� �M���F� Βu�.�q�f-^5LlU(lMR�BZ���K�,�m�sT#5�d���Z��������tiiX�:x�D��GЕ��}��ʡ��c�Jٵk��5 ����	@(Y�(�p�89ò{���im�����O˲�˔:Ŏ��+������r�_̸��BzdIGas ��*�I��� 왔%���{}����ac@O?#�w�#D$[�)W�U�9�O�A��`��O�@��3��n�j�-���`ri�������ڎ"�4	��w�f.Q�C�`�6 ������{�z�Yh昍H�n�l�������� or%U!���L�;d���Mj�,GlU
fQ�mo��g&g���k%���^��aQ�@	H�<�ȼ �4e��h��#(��C�f6�(��T�������(کl�Wd���L�'�����@�jx�X�}p�1���!:�Y;�k-8�9����1�@rX���N �8*oB��d��B@i`�9B���t�mw'���iZ��C�ÿ�g�B3�'-y�d�H���2 �lP>ô|EU����v�?���6�)�̤�Ӄ J�5 ����k#8iim�G�OvlߦY��1�,
?�7�rfO��'>+�4[gʧ���5��Uơ0b�,jQ����r��r�5pt1[s������24�IXl��3��]����ጌ��V׍w�%5-�djp�w��eL&� )���Y[���9~&¯Y�y#�QCWΎ�k��%�JORfp�m(ڳ\��wɖ���T܄��.ykS"�.�a2Ji�9� e���X����՜_Zxe��Q�2���y�Ƞ��d̘��)���IW��"��_0Z�V�F](���3�� �5�C����7�H���<�����`V�³�0�Bp:5�$, 5dL�i�yq�Ұ6�\,H���f�wk��^���l����/(���ٯ�ܮ�Ո����dƘ3��>�z1ZLFs0�~e���r^:�*�2Sȝ���+ʫ3��VoT�W�I}냕�kvj�mx�-��QN�e��0��E$�Lɢ�u�`1�!VPbN�A�D;%�-���6p�%`��C��R�{9r[gh�#��=po�,#�1��Aȵj�p���M���⭞��˖Iݚ{��Y�S��4�P�����J��oÞ�u�}B^;[����*~}ʹ��m.9`Ҕ��n��^L{���O���3���4lV>�D2nB_��X�8�u�̻}=0Ń}�1[���	f␻�Q %ϟ��|X�Ĺl�jH�g��$t�ҩ�
&kc��@j���a� ��v��ڰ��>��]��=��q�����1�a��.H�Wޡ���a��wd���Y�:Ȃ�6�m���$@R���R=~��:H�?I%��'� ���XB�A��Z?�<�d�`E�7�tn8Z�
Y�8�lM���]X�����%%��
dF�$�����٪E��o��[�3�s������4s��T�_tL�.lW�k�AS��9o�5��̙���`�������P�o�eX���.='��,0�W#>�r�j�5|�]?RcyX��������n
�e�v�F$����ēRc��#СRd�����e����D�: (�ymj\�N=H,�����r�-wt5��)��̆��� E� =v�����X�*�
~t���1�ܢ�9P~�
o�T��E�������Z o�F�����d�hS��S�E�_�!�W���T2Ń�*�ԁ@�Y�6�o���[TpMC�%�����F�R룶�ʺ��93���z�����yޯ�I�'��o�]�}�y ���_�X��#�H��"C��r�hRN����>���O�\ƢbuK@��� `U%R%$������6@ׄtuF�kZ���cT ��$�B��g�Lt]*N����1�џ��$����+K�l2�vW��|��*��lBv�$��zR+~<���e,X�E��6Z�T@�z���(�NZ�X4�+�'�F����(hH9�#oaZ���7P=#�[`E��?��=� �:YBOrv���8�қ5K�x��)9���L����؝m�ֶd��Ҷf���p�,ת5��@Y�k�{��˾�4 �3e��4��׳o���`1V�2e&����:?gi��U��$�3��r�ڐ�H72�(/Vj�Q~�x>�e�-�������W����d�a]PŇ��tA)0�̒%���?.����5/�) ��y��O#{�nB��˦D�=�z�����;ZM`b�,X��F��
�df<_-K@���(.�U�"�����,玃�R�T�0
r���}�����u���	�OU�O�s9�a�R`��#©-(��y��I�?x�8����W�����\�@��0���ƒ��ܡa�8�-|�L����ⷜ5��A�*eP�d�,Ƚ�g����sW������<�=�G��5���މ��@X��,�UL��a���BE|nxn{��t���`�:�'_�G���b��wi���^,fdSNȾ�&;�֬
�j�*>��rz�D�i������,Ċ0��p�a�Y�=A^,/\jdw1[ȱ�!	��(�����N�jY|�~�B���fV�ï����{�24��B���igpg�$d���e��?�L^ւ3p�H���)h^d�6h�n��S��֦�`I�'0���������:�>E�Hީ첟���(���I�wGP�m]&���?\�tM��E�v���Xq5���3�����,[ձ�J�OCkދI�wrL��B��E��� 6�5l�i[�Jj��@]����E��/��Yf��eӚ?����}���o,�Ȯ��-C��.*&ć�k�<�Ր�i5��u,��jժ���'�P�`f@��ٙrL�wp�/_�J�l6.��5� �b&#:�{�o�z� �y�G֤�K1�>$0N�Y"����|�@ٮ�C['��'`�B�AV|�J&Z���\FU�ܑ.���%���z��Q�0���l=�I34�*�0Z7Hf���g<q83�E�v2��?6É$��']���X����mq���j��1�v1N��M��Cfo"��
m\K%���giw��n.� �+����\/���!���{��}v'��m��f�z��7H�Y�9g{�r���� @[Z:�"�f��ƀ�T��e[� I^
��]�'٩>.��η��}�`AS�)ܽ��]��Aٲe���8U���"j݋�~��g�e�_S�q#" H����z�oO_�=zD����/X�������ݷ��-P�=�PLXC��%J�`�Fzs<i��m?s�LĐ������Y���´�:N!� �۴\NB�D`�V0�1
P:0�X% 	kC%����
�	����pľ�	���z(���.��㚚���WI�F��
���f��*�Ī��#�ٓ���	��ٖ#s�w��q��l���n��p�_���<Pɤ�3��E˟���}I�X�eI�N���h��@j&��(�^(��	O��&���
����ÜX���\_��0wrB����{g	ï�oA�m���`��s��ƫ�z�X�Bz1��q�nov����Z����5��c��\30��>����rϡp�Xg��e0''�k��*�m���<�/Y�,���Jiu�
Ml~���/��?(o����!����%(A�� ���b��{B��]Ę��k�Dn ������ƴ2=��ɓ'�7^���N�����(��
+���BG��Qp�xIV8��G���ݫdsGH�9�\3���������g��Q���Z�4,;PX���2���r����+�1�����wAuR@(yব��ODX��kknح廑���
SȜe����u��i���Iʱ�Q�,KS��8�T���1��噧���NE��FxR�4zS�T,y�^�A(���}��wrE|��Z��~�8!0f�Ekc�p:c�(��S!�� U��7_��,Y����;�7�����T�q�X�U�]������3`
��b`�M ��e�ĥ���F�c�T��������h��.�T�53�B��;%]\��
>���>u�}r�{-"��/�#@�LFm�+�X�'X�Ȓ�O����)3�X?��k���A��@��$#t۪�ɯ��]Z���Vٔ�<�G���P�*Rm-��Cݲg�+��K��m5jTݰc#b)z0/h�f�5�� 2uN���;� }}�H�H��>�~�SA���QC=J}��� ���z(�u��ltw�ݪ;�7��x�a��T�3�t!E�ow[sٜI�F���i��.h;M��M']ںJ�u��x���_�N(���ͤ�H <$�5]l��{۫�,v*b;+XB
֛x��]=H��}] �7	~�]�?DK�}��zh@�<6X+�uI׹Y����������	�&k\C�����9^1���p�ٮ�*�T��1��Jy��ay�=C{��S1� �;3��6&+4��|���|���׆��l�w�~C^��W��l��6Y��/�X� @���&Qv�-p^_����`�^�&�0as��<`4s�{鄃���jRM���!`b��f�]C�{e����̷-��F����]�A��Cr�ٿDu�C����'z�_��!�֬��_��� p&f &����h7�m�P`:����<ݫ̂۵�Y��Z:�y�[�Y���N����?�����)�(��q�78��6���m��~�^��OM�[c�>���- Pa��'~J�;c�s�e���Y~�����X��c
�j# Idr?w��{� ,M��������K��8f|�6��)$Q���󰦍��d��T~��8��~7�:�c�������/0喝���|Q�
i`e���Hc������!9��E�!��:KI�V��#�U MNvKd�-F&��]>I��ȃ�V��p�z��ܡ����������U�^�:��#Z�8d:N����<qI5�w< *���%��z�>s�Kw*�A��};��ޒ�9V���e7/�x�������hL�׾��J��7$��(h��as���P��J�I11zD�O���Ki΀�j|�Q���i�]{B�ŵЬ���p���n�jT�V����Sxf$��e�_A����x\Sa�?����s'���au��`�P  'r�H�F+�����057�Ħ���%g��&�oA��㨂>)7�	� 2'� H�!n-N+�|jdJ�PT1���!kv�au��p�̡�|6�J�K��E�v'��o��-(�jTˀ�p}y[K+��,]�U	r�zT@��c��3��dGv-7�+f�5 U�8s�ٽ�=�$8L1�rB��ke� 	C����=��d�V���r(�5��Ɉ_�G���K"`dB�0�����&q0 ܖ�ZUhyV%�|F�dm���V����m���$������%���Ua<�![8�����;���>��a2�+ehhP.�����&��/��c�)%�$��Q2�z��ۜ`�n2: ��Pb�*^.3UAt�<���e�^���,��nwZ~]Y+�%�ǲo9�Eo-�Տʾ���c�k�dݖ�r��Zʄ£��'#�z��)�֮�6V�J�34;
7�1�KL��3<(8Z�+����-��W� �6�G��@���~�>��U�x�9kb�	G�J�/��t�n��@�b4'_�s7=y��c�Gi:d�9�1JY�.�:V��V���������0��<~��3�]Ziw��޼�w��׽���@�$$��ABH��ϗ�$_B(!�-�f�����z���ծz���H�?�9���F��-F�+��=������y�+��$��<�q��URX}��w��Ʌ�
V��|��r���	A԰UW�ȭ7�$�MF��jjAh�怦�/>B��R�a��x�J{EO�� ����'.X�:b"X�J3?>Ȁ��i=�gkW��!J��l��ɨ�h�Lء���c ̠�=1��Ѱ*�)S�� OjK��Z*��rON�-�R��=�����{Z��S��/>�����1�SY�\(\�t�o&���o�$#91�%m�Դ�q��5p��ҷ����A0�/���5Y�=ݴ{`� �E�9���M-5�!�|#On*��(6��m�~�9��I˲erϫ�ATC�af#�0��v�!)�us��H�0�	���}RF(-S��F����2<�����݃��R����:�X[Le��{�lO#c�$8T�҉$u�ܭ���m啩Y� HVQI�X�h9��G��۴��I�4x�`Q��*֦U�^��޾ud��}��P�G$��8��V���KI�P߬��ri�>�<k��6�2�-/�������'��  u�*hn� ��P�C H<q<�@�d5�M�0R Mf�s�t�`�t��\���%�}�X�'xֿ+�,��]9�7iJ��9Ѭ���&�$���P�I���$Vx�TV=#�}~�Y�g��j2XT`?Ձ'Vp��e�?��S"]0��/�f
A(4_N�0Hg3�w\��{F�1���𣲦|�ةiB&��2�=p� '�4�O�p*�8���~P&+xZ}�G�N����0�T���+D�٪��)�'�d=�~CE�:�����計��w�{:�o�jp��J(2-�BzC�ԁ����uP�K�Y��
�q���| �5�<i����ۂ��?�N�vG�44.U�3�T57����rQY�q��@ϓ�n468�=�1<\�}�(X�^�/�g�
o@�n��G���X��G���䦛n��:�80�{��
܄��$=�z���ȵ��gZw�"��p�Ƈץ��t��4��e�Z+jn�r�h~#Bf�I ����s�����M`��]ȯ��:��������_�0��կ��Ÿ���] ��(X��!�6�zR�%e����m�իZj�;��������8ӟƔ�ǘC|�2�`�T���r�I���������ZE��ݽXC�p#l^�&�	�%m��C�7h�w�ZhJ �̖R��Ҥ �``��Rbwp����5�X�Jj��\�&Ǜb�G���=8�i*�_�#��#���kOu�ӯ�2�_!@���⪑�E�r���~�E�z$�i���l�@�N�s���D���-��ʪ~�������:#M��d��o�~��	)_�ڴEؐ��2���Q�Q c, N�~i��� &���>p^~��R�h6 ��7����Eo2�
$�� +��մ���©��;�y��t�C`D)�E�1Q��Zۀi���7#�Đ61� w��r�:�K���CCC����.��ӗc,�E@-
�7����p�-�ۅ����K�����A��C;pD=�T�~IĈ:�G�!н���(�k*q�(s��\)z436o�t���f�&���P��
��3���̰M���ch�p���<=���*��[��--���\�v1S��a�Z��hX�xɺ��U�р�z��*���������ڱSn��jY��0K��q>�0�r�(x��apD��u
� K��!߅M����@S4�����7&���(���K� /���_d`pk
ίtPUЦ ���&�����*�+�Z��WH�	F+"ʉ�q��V[:����Π��ϵ���߸}�Pe�R���$w�����9B��8��d�PUѷҚjC;����W'�fX=�M��y SQ^�)���P������Ř`�3�ٺ5�5M� x�OӪ�%�X�F�d��1 �� �mHH� �#�F�o����.�F0�L�(��G͒\]��\.׮�Sqû�k^��{�'p^z���N��(� �j�C�7+�IS�VD�$�K�0��0�̑L�b��Д���M_�'�%���>h�DΜۏ'ߔ���G3��t�$�qCTq�2p_���|P�GӒ������2o��7���l &-')��@�#8�� ��P�S�N�Y��A��n���$��%+jN�5�,�# l�}ȋ��S��� \�Q�<v��i�hJЦp"*��#r��0��WJ���А�u{qW�)��-�����1)�ںAe�kl�1�Þ��\�ދM�-���f�
���Y"��"r����S��p��~���0bF��9��~�����*sɺ�VY���|��`�>���_����������C�q����xR�O�	'^lTZsPW�Y®m�?�8�d�{*����Ax,����K+��ĪלM/�y��L�q������� ����H���&�϶��S��A�����R���?�����J�9F�O|���wf�i7U��{^-	8�
���;[���=����i=ߦ�)�
�~+R
��|Eʗ�/N_5����õ��&��TpT.�A�p)��o����%�����e>Sʈ)��*5F�������#:���>L[�\'+���#U��Jg]��/���@��'��� �j��J�ʗ4}YR��?q��R���BN�q%\Dߞ�(50/<F�LC��HJ���M��ƛj%D��L/�/����_�����Rd�:�s��W0�Ai�i�$"�7ͻfS�׀?bhyV�ȩNmz� ,aF�Y���K\�9����x�=y�4�ҨJF�eF+ОA��Q�8�][d�}�k�' {��^)��kTʧy�4G�&���L�RO��:�J���D�?���F329?���PH��_���	=&��jDq4��I�s�B�D���9tTUJ�ќ�|c���\�lebN�=�1��b��b�t����5:���q���񾎹�FЇ;�5y��S�R��C�����I��x�)J�h*�5��B9�q��`��8A�w!��Q�6"���2�áeʤx��7iw��>K�Ɋ0�d���}�7��g;�	Sp��������T;�M�����c/�:2q/�)�7��"�V4��-7�#�p�|�K_����,��o�18|��L����L8����R�ˉ��~��
�r�����d���'B��,����K��o��K�kks�������C�C�����:z�x���Y ��B'��@���6�S9�:s�U&�ΰ���p;��:�P�\��S�a�fj"�����w�S_�}[%�KZ�u��#�7(ͭ�@��,�E�J�xv����0*�Bf
���hX��~-&ԥo�aO�|�y�V����5�	�v���X�G���I�35�i�2y3��خ�,u�L��r�>̓Ÿ�G����@B�oZ'��9
Pf8HȪ�VK�u�$��6�f$�袻�k� �#c��D�9!eU��՗s�r/$ ����K%���S>58y�t,�h�1����̈́�gV�)U��.	���eڤ�:�p���4�p�K}�"q�b"=���g�)��O��\�;����%�~�vP��#@�!~ -s)2l�E�d�L��򊟈�0�����Ҽ��V����|�u�4P�׋h���?��5�������A09��<u?��]��d������A�o�B���E�&���r����{]�l^Y!��q������j�N~y�'�~D��W����ah I�J�F�
#�h�i��~6��RO��6'a���?i�0���&����_QS�AD$)%�v3��/���Yf���4�>a��1��Yv~
��a����KK/�c�(���#� �T�0�"'��R���������#�E��,Y�iޱvE��s�&�{mF>���e{�+eba��Tf�I.�C&�.�+2�eT$�JvL� ��&�����
����� �f.j��~�qӄ<u|���@�Cօ	�x@9�^�4 n^u�K�$��`�j�v#����.X*�ӕ^0Q�r����OJ��^�@
�nSV	�F��ڣ��<�2\7 �	^�#��5M�ͣ�\Ee�l & ��	4J� ,G��-����w��<���F��C.�
�����?!����?+1m�g�hlu�����&����,ftV��6�t9�:,7{�Ѫ���A���,�>�qZ��ʙ�Ҭ�� �����C�(�M�=A��O�ɟ��Y��D9b�䘴�&p2W�J\|�}H΂��t�_����r��F���Q5�|�_=|@%��yr%J�DbTT�$�d�xz�@�j?Un�F�-�ǓvTJ���"�S�쿽�}��gu_�8f�{Ă+�s-C���u���8A�Σ��3Q`;� & �FR��g ��R�15c�;��Dǰt��"[�K���AAS�����	�2������R� ���.��{i@�Y�$����USsރs� �ܞ����R�*8|�w�+}1��:�'c �uvu�Gt|sV>E�$G�G�i4>j�L�*\�>���r{�|�k_��^�-K�5H�5I|y������g>�i9s.���I�R���P3b�-��zf(0�}Yi��wli7�����Z{�#�*��;��H`rG}�e�}	��!�	ˤką��H����#4IL�F�����mΧ�+�3L��m�#�`l��$��I<Њߑ�^�.��/DM�Y�y3j���&9U�LTF�a�p{<I�.y:��@:g�Zљ��w�����F�9�G���W��KS]��_��n�������[6"�Ƥ�sD���ii�/��"�i��I"�0}p�S�n�䂖c<۸�)LO�2��o�i�oN�������L����H;^kad��2���I�	L��n��;&�bn8:3O�{���@`�!�V�j���4��׻b����&�F��v$�k>4�#Њ�)���/�8�Й�+ajo^�$��!D���D�9?s�tE�	�148 �����2���	L#$C�9���T�=��V}NkЃ܏��T^��I��z�� Rǵ�]�ݶ��3tG�Z�S'OHg�y�[� ˗�@���O�*A�{L��9�<��N�рW��N7
�*����Z�����R ��d��^dc`�!#�<t�}�T�S%sp�ş��O�1`��F��s2�Ն��Yأ�=I��*ߡ+�L��Ȼ����x:7h'Y�[SD'�	Bb\�ey@捞Bcױ^9�>�4M���w�� ����?���*���N%Æ��FT�_�/-���]���Q���� 8�f�~f��뮜���3bW�=��b:����6X��ɓ��Eu1Y�cj�D/I�2�O���5��Ⰻ/��46�#H�ǭ*gq�l���d����!��W>V�=�A%Шm��՛6ʑgwK�h|S1V.�2�(�F���ɽ��*�Z�����ܛDNt�e�(}��/7���v�\n��_*J����g.Ȫ�S��:ա�-Eа�����뮕M��R�������y8a��c��RQ��=9	���)��7`ݕ���3]��R��t�vό�`�����gF.�0	�6�V�h"�9�f��'�ك8��c�곆(�d>P�=Ӿbu�o�
��-5�>��Q�0���.��h"`"���,�i�������yM&��J�Y���mn0b*�;�0�T�7�[�k���ݑX��Z}�8WHA�����F�b`�=^��9���?���׹�ƈ�`Z�9���lP�ʠS'}N/�~�..��VQ�����D"z����2+��Ȟg��/rM�
� �����$���;NY�b�l�z T��I����l�[�~3�8ӻ0na��i$�rي���(K�p�+*)���r��)?[���b�h�-,LQf�j/R'A��LT>}�{�E���M�f�~��_[;j��[$���S�:N��Fes�Q�P�s������ã����^���i~��H�[��r$�P�X?�_��N��\S��׃�� T�����1f����ў��u�]m��ϋz<�a��� �n��|�=�p�������vG�.��f=��k��>��M�uuw ���2S�D��
W��ytt �)��,܀�����ٽ�H��S^�B{?��l*7��W#�Ma7�3K���T\�(ޜ�=�_���e��A����2�N�\�s��ֵ���6ܓ��j�J�*J�c��k!���R6�*��K�Ď��l�ߋ0��M� %t�����؁ܐ���1�䔶;���&��x`.a�J#��--+UC@����V���%]���Fny���#?����*��D�M2��l=Mp\�sAs耦�S�9 ~����0�Q��BG���c?��a��3�)���_1�����r��O��}5�0}��}�g�\~=����}�C�<��7�i3
M$P*��H��X�T?�=�/߄��^�R�F9���$�8�OQt�5g^�����QYz��j��C�5CJ����D��'QU\~�9�-�� &<,K�'1�T�˨C7��h:S?[|�&{Q�j7"�`�fIm5�̷:�&B��J	|��}�rq��.��VɃk��dT����,�wE�Q?;�(5/)��q(�~����B�,/���zy�OH�o$é&�m8�{�
�Q0����E�}ǫ��8���e��d򢴕�6�����d�/��P�U�TT)ĥ�멺S\�o�UKƌ&�}<�N)�������?��9�'�ߜC�0����K.a8�.�t���0Y����k�M:�>"'����;� ?qTn�PB8����#C��F�Oy�G�A����u���Ң1Rφ��ǉr�-��:�y2�N�J�^2���
ʔ@4�N�Ù���O)��ǚ�QM�w�����5��1��$�׌vj�p^��;�גb���&2�{��j�sp t	:�3G�!�l�(�fW�2'��k��M�񷶾��<��d�c?���~.����{��2Z�	Zf�d�U�>�	��j��	Q˂��In3��%_���n��ǆl�!�8�N#��x�B�����WE�]`t�#,��G^ �M���^)n�A��<>��%l�+�ј���/�����u�Xb��v�!�̹��(-���")v'�����h��Cp<w�[�Pٻ��3���`h�k��Je
C��]���p�И��pC�QQ7*�ZEEEn��)������CkVR*�'z%9���3)W1��[(�m���@#�&T3����\qM�0G��8?҄�����R����奓��A�WC�׻�AV�X�`��n�ϫ+�^�~*Q�t�w���N�w�#KW������ثr5����� _���b� E�d�(�#ਉ��`\���ы�J�@ʌq���9prD������JKL�;��C1��ʛTi3�7������0���CK��#9��ȴ�¦p?�p���Z�س��|�-�)�ӭ�r>G��a���	��lk��}�;��9��ɫ~�^���U���2w=��G�#�n̗Wx$��g�L{[�����f�1������GH1����L�HP 
sO�XK��d1mL���,*�O�UW�n���#cw��3�N�}*�E��[������91�����z��H�Gz�Z��������s��X\.-- E�D�O���Ct�,&��2I�I%�F� ��e��!0a"i��a�y��,��}�t�-oV�#�q@�+?(��Q�Wv�7�]**�Y��a�)/���^%8E�HO�� ;j'��}J�A8���bԧ��Q�c\����gn�gN:WМ3_3��x�s�֝��v���O��L�;͹a�F5=����㧲+� ҭ3S�w=���,�0�H���KO��H{e������O5�(�*qa��=��Y"��8,`�������<`��G/���U���0�L��|2�J)i���)���ڵ�����x�_��P@J��(�q�[�Y{�Jy�m��|�oр+q��{CH�@0��zi���Q����əS��*��L�	RL|��/U��*B����
�Q�`��ϸd�}^q�-�g_3���X/��ߙ�Xb?��o	���zV���0�ں�Ҟ"A�;���y���{���H}ci�#�MɁ�^���Q��X�pƒ	vu-��n�&�� N��KL �4ŭY�\��,P/���4��J���hS%�$ClM@�
X7n��V�(�("H���qe`z�}T.�+M����\T�G�"����m��Q�'��4>ɼ;�Mc]1D.ZpQ����l��- B�Rpp�FaT���Q��ȗ�֭�_H��S�?�B3�)@�� �FG��©�Z���b�y�Ż�l���u�w��C�i����>A�����du|�*t퇫��Wgl/�;65������ǎɓ{�$ ��φ�#�Wnh)ǧB����RE��{I�����G\�,�(�� �9��[�p$A��Ge߁��ē�+��=��W>�g�Lz�(�}B���	���#�7�|��p��le���oGH�����'��~ﻊ�p�������뤬�L�kQ)(Ƽʬ�^�����.���H��"Ij�������4����h@q1 ��I{�'S^0��i��H�� %^�ڛr�uEH%S	n�Y�@L�g.7��K����"8�E+c�y��`2e�	��M��Q�Zp|�)=�fk��>=	�RT�3�jΟ'~�K�Oݗ\w�>�CnY��N��ӟN	���������� �^Y��V�Tޠ�h3ZP3x�ߖ[9�K<��y����,yy"҂Ų4T���;&���%�,q˂J�Yx%��Aq��W/��7րw�/���U�PCM��[R.�k}R4����2�6�8���VK#R��
m�9{������r.�ʯ~�|\�a� �^�yL��+Jh$�Y��}�|�B��O��� �k8�B�A�;��i���G- �����#�e�����F8��� M!�|�J��'��!Ӳ��H�0��O秴�A�`DA�:�� �h����ح�tѺ(��(��θ�;�FT����]/�ɘ�k��$��,/�w��\��/R�t'��jT���fEE�gL�x�ҧ�Ў䘡=^<�I�x�<�g���(�ys��h����d�P��YJдy�uʧ�.�
ө��%Ҽ�e���:��� ���_��r3��Y�J{�y�4�{�U�fk˭}�p�~�����J��vq����Z��ii�V���*�����&k��ڥ��N��&����S/6,�������n����+����m=��O#��+]V��h.l�������q}�{~a�~ �0�Sm�������\0|v2�[�s~�,������*[�QRg
�cnW��߃IJ���f���8x;*�е
^�V��IF@Fm��0��D�8��iXd�koA��U���C��vQ/�cM.¡�-w/��/������]�\�q�z%	 ��2�|�1f ��-`6G�zjU�t��5U��Q�z����dl���qJn��*��uo��m�#��d�@�b+^����>���E�W�Ô�L�ǹs0������6�'l�!�7���Q-W�����SU�FR&;Zq������r)<�2���`�QP�5����N�,ʄ�t!�>
t�˭�r陉�0�L
UY�nhh8�4�)�yhgx�T=��rލS��)w\h*�/͋�+b��̛r(y��/c퍤?���vL����&*�-4$N;�w�*.�I��= $L{�K^c�8e��o����?e3��gI�G�#;�d'x���C��&�MG�O�L��Y��(��t�x�?�_��5�)CL`����YH@ͺ�	�F�n���r}K ��9�Y��3�Ԁ~���^F3'u����Lj�ˡ�2z��M1����>R3o_���:��d-�l*�|��K��]�����2�J�`H���d) U	�-����-+�������qs�fZ��s$��%%%�F(*Q Oo҈�����A��Ly�f��Wtfi/�:)Gz�/.d�xr+~v�\�+�%ndt��(�Ԯ��􂲛Иy����T7��^����� Y�|rnZEX_�pT	�|
��XO�i�_�m ��U���r�6��'kL@S8�QhP�׋��^��?0��~s&?�mm�w�ౢ&x�;Մr	�=�֧�Z�* sL�Gp�U�冦A��?Y��;,nDn��=�^�-��r6ĵ<�!`���W��)@c���
Y�q�476��I�L̓nW����Bs�O�3w����m_�N�d���0~%��5#S%��h��1�a�G�q�Шm�eOG@^Io��y��髯��k�����6� x� X2	s�9�:$?z�U���W�9F �5�i��>0��痽������;��z�2M�$u�a�,++�`N^m�E	Ws��/���x�j��_Q�=JkB�����+�.F22Z,�>�G�748�:zl���\� ��nl��KZ�&}�����t�ܐ�;3�����ehF+)�H�r�8a"�P,�C�B��	�ܓ^��;fO�Gk!(z��	�ƫ ��zN�׃�RS�Rt��v�T�)Б����|�m�]�wߋr��O~��W)ԑ�vT�r��&�!��f�?x��jt�e+|tV�4+m���n�������	�`!A���8*���)��쑿������&��A.��ۥ��a>ͬL�jY=��re���}�-[6I,-����r�kL>�ݮ)����q�+���n�kr��L��3i���e�*�h��*K�//�/�֪Ee{TyzԲ���n�"1O{o�
���S��;�1��!]@M_Vu���6'wq�{�k�z�5Ls��WV�Z������˞����d&
'6�d1'�Z��'ۆ�?9&��oY$Kꭾ&��5	*��8)N��w��E�#����ޥ�����4�u�-�2��12)�0N�ēK䉩�["�5�e \"�^�V��YP�ٓ�?���8m����������h	2�DĎ�:n/���0�-�@O�(��%�w�Z�w#���z��d������{��e@Z�w�}�$�L��)�25������L�(ʄ��0
 �^ ���x��#r��F|�W�5�ߪ����,�Ap����eh�(8#;�*�-Af��y˃rۭ7B��&|����L���tT����OS	#���" ���kG?6o�OV�Z"C�5�ͩ����!���q�CD8�q�&�E�IXͳi11�w�,]����sG-%}���tf��ʋ�Kv]����,i,�}���STʨ�>|�������������87`�7� ����e�yc�?��;�~���
�}0�=�B�\� �\�{R)��5K���8 ��BHp�HD~�/$��&����_J	 K�ƈ_P*G����ť���2;�$��S�|��\)�f~��R�:�g�7���さ�_�c�#Ȇ�����Q��I���AG���M�/���%����̂%c��c8�),`�m��A-���O�s��
�1$e2͕P�w߽�7�^>�ῐ����ǯm���.<�b9j��/s���@��7~�Z�L�J��6]���k� i�,x��pL��;,իo����TW�)
�x���LG߶L��(J�����75*�[1�ȩbt� �-�;����K�{�G��DvVʦkWʵw�.?)n�21+��ۤ�.1�N�x݃��[l'�����Z �:����n�0MO[�m���;�����p���Y娋��PvыS8�Ik�<Ͻ����ݵ�~0�'o��)�ͯ����g�G��_�,m�D5""��"^�y�s:���y�t;�J{Tkǰ<��yi(�y��F��@��n�J�I,4�ӝC��G��A�U��	^�$~���@T��Tf(�T=݃�j�iT;pZO���d*�~�ؠa��F��ɲ��L���x4 ��,��I���E��Z�!�A�Š	�� 	��4Ft$J==T$��}*N>E�;('j�/�l�)ա�ʜL4�y������W�	�/"ϒ	�*x"�×�Y��>qj3�6�!��
# ��i��@v��w��B9�[��d�N�ׅ}�F�s��`^��$_-p���h����_���
�4.iR�Բ8Q���S�7�<Z4&�c�ؼ��n��W<�+$���H[o������p���d,�m�n��ͩ8��|���� ��*���<��`��P !���w~���&��J?��8�s�1( {�&f���m٢Z����HeE�jc��y=$x����HR�Em�~��pR�V����ߑ��R��!),_�/���ayQ�����,��^|��4�dV��w���{�{>���w��`�9�ר���N� >�!��<`��+�2}�2PX7V�R��`�$�#�����eyS�,����������>����ؖ���-������|� q��'�����:��6ӌ��O��5��"qۖ��I��+����k,������9�
A�۷$\:;;�o�ߗ�x�`��N�F?S�����B��r8�P�O159ɱ��	��=�Q�7�\�NE�'!+ا $ r ���)a�&�����	)9��n$�+��734��]�>��qEsuqF����\+��ݢ4E�������Qt�y�����i�^���2� �v�)1��@���*��V)��V�r��.�z��*3��D�4!~��o�^����r�;�M��.���T����j&�L�2����u0�a�s����E.�a���".�}�����Ð^9�8�]�1~�z����K�=�0��+
0q���� Z�WԢ �5��{�,�5��P\�ܕ�]3�zp�,�6��~��ť�5$g��y�'�T��t�ʺ�����:	&��PWևMr�!*�ݻ�����M���t+����/}�k���������x�U�Yx�:|Y#]g�1�ZEu�yi�Ӭv�eZYnjeNߞ�a�w�WJa�cd�>��<�{W���ɻ4^�v_���QD���ˏ��`� �Ҏ�� ��ߊ�,�S����o����}C��gEpG��l�C�`䋗��"�� D�����9W�'�sO�Po�T��]��8Ͳ�d
�C�.HMqX<%�tEMC�g��RqLS: i�AoS8�)h���A���RD~�����W�����Qtp`�bN��C�7#�:�wQ�ho�&�A)�䔘�!D�e򵠙�x�#C1�l*���ɗ Rt=���`:��]�}���֩���hO �t(5�.
n��d)�W�C�auǃ^��g�	�[Ag��&D"�h,����+�� �hD�"N9B�fe��� ���N�߇~��ɛ��JY�kh�`���ө�3�P~�ԡ� S g,cj�دZcU g:��
@�:�Ԓ*=�3���n �� e��\� �n�k�h��*��զ�I���0�~8׷i?N¿�,,j�Xq��|Ƴ͞Կs��N���޽�w��{���/����{o�����>��h��1���a�<��w;���k�l��|]z�ȶ���\�rJ�4&m�A�e ��`M �I�lYS5Im��.[WU���ݲ���:�!�@N\��JP�5��WA�c���o���\�Nj�0�6:2�f{�����̳d��]Ȩ��QDO�ĲV�_	Gp�����5�K�rN{%�HHt<>mx����7��,��3�-�gn�B�aJ��d��$���z��`�&`d1�k�����:-�{�[�c�#:K��@1hJ������\��.+���Q.������i��BcE��hWӣHٞ�ꍹ�?\,��#*�W�������J�p<��*%J�P��^'�:b���b�K)8��b�G��O����#.郆��0�D��s�1���7D�Z����ƆwW���x����ehd2!���R?��j�q�y-�� ��r�3�G8�'A�U�|�<�.�t�F5�0���$������{O�j^(TF��l4?�-Q�S�[͂�5],Jhf .�u�r<�	�ü:��	)��,���e����^�{r:<8���Bo��,�A����o)*W���u���X~���ھL����}���������gR�d�����ׇ�{����rw���׊��	x���fe��A�7��>�L�{�J�"׭6�=;��M�uJ�I ��"D��$!��3@.�)� &'�&�8������}'o��Ga�n�)�M&:�*�'cS,�_!�*�ze�� �u�}�ky���j �j���CX�+˥l�:)Z�A��T5�n�%���T8�kQ��4ɣ?�E�Atxd*&�I��� �O������=��WV���%k��w�X��o�ING|J���� )J(��$�\ې�;6�JM�"y�7屳�H����������P�V�5��X�^���D�h/��$�<�r�3a#5�fnK�~��L`]q�t$�qd
} � �?kS[�>[p"� �}�d�_���J�^��� �4��4�73��w&���{�� �~�6�pʹb�F�}?�p.Q��ޤ	��S����LC1kO�	��R������9蒳���/�`9*���d���5�"�y��E遈Wʚo��:���&�[�C�8�AC5�V�dw��|���ٳym*y\|�M��}��3�ÃUc=/��i:k�f�<���K9�0�����e��iֺ���(�]6��A���Qs��?T'Î��I��kW�%}���[��LV��S�Hݧ�ߴ&N����]R+�n���G"#]ꔞ��*¦�I�MN��T5X7n�V��a�� 	@��%{���r��J+��z��/�&,$&MJ7k�ږ�w+�U�\$=��>"�B��]%�5�c���hz����@�_QJ�!i�I.��K���*�v����.kAk�ܪڠ���oʷȍ_��$���ǲ�����6�#?����t��w_'��j%�C0 7R��&eI��iw��cM�8pD��>��������F+	'�/�"F��9�T�C��h��C�R�A[EP �$��^��Ԙ[�ߋ{���)��ajޚ�Z*K�f�D��t��d`WO�����z���Q�J=���T��
���ү'�g��V��{�,����2b2�:y�$�{8��7W���o:�.hZ�DGG۵�B�D�w��N�l���b:���j�ʋ��n��f�7����8�%���,�Ҵ���"�!�|���E��~.�7�r-4�0B�d��bw�H���;3/U��;�2ջ�a� %�$W��Fa�����*\�_�M��:"k�6pi�`� ����U\�=�w���L��&���e�����x�"8��ʷ~yHڇ�J`��O�'|/N��&Fg2R�ڃ�K�h8�
T#��I��'����c�~\���m� �K��xP��>}���'e��#�M��n)�/<V RV�R��ɗSNm��9ݚ�1n����S�E�&�I�Lp�p^N/��t�d��Í�p���|�\��Zk}��B2Lo�æД��T��ؐ�˸�q/j.���$�����U2���%�^�m�0���j��W�R��+8�ꅙzq��[������~׭����];_�?�D�������n�f�E��3WWr֔{�0�Ls�ӗO�S�q�##��NVYP�&= �`�����G�x�����>�tXxc��:���ҧJ�jH�Ѕ/��f���Zr�De���8�1���f�yh��s&Y�u4�*2k�Z9�6d1E����3���ȡ-/�w�����'g���<�,�KZ������G��j�>��:�'}�;��W��%��2É�	CЀ���H��sȱPb��K����}O���	'�ߕP�:C�Đ7�H,)Dy�F9��r����%-�rp�Ap}Edٖ��3�/��/�v:�.��#C��E��H�C��� c9�|m��sF���L�D�Vixd���7"O�~���h�GQ}o,8�V����6RD%u�J�4}�����ˤ���Ky��d�����ۤh����q��f{;�%	���
��U�t�톪����_��t��.�kh8����"�p)u�`�ۊD��@噵a��9O�N{���l�y�<`�����jͺ��T�3�x2SQ�>�������5��H�PT�*�U�\Μ]d��&-�4�]W�~%3$<���g6ȽމWF0F�� ����\QCJ�j��ƍ���}2d� \!4�[�R �T- �J�Љm""7�"�Yyv��+�A��9���n��t����i̤��a�|��=a���w*d��J��K�N�qO��pjg席R6�S��\ޜ�F8kz ���ġ"��ߗ��B�=*i�[֮��?0E�a͍r����d�=F_�,e&���jfB�lϙ��3�9I��/�Vz�T�������bʈL�d����3�g�}�M"��~�H�$�[ڮ��-�{+i�cd���K�Jk�x����R�~��p �`[��Ǚ̇�ܻ���?�qO��ܛ�=w�uoϫ��R:d����#�����3��r�� ³umK�q���)�~�^�.=�T�� zE9�b�<�Wi*���E�N�i�ĉ�X�MR
�B�o�_�L�o5�(�dl��:���&��69��s�`�pRy�@�7�~��i��V�F��4�i>>
T�i�kp�^�"4�A8]sn�݌��|�E�Qet��d{�=�[�!�xW?j��L�5cdnV��q]��Q'2�aG�GA��j��B'����2r��(Ӵ���ʍ7�Uh�z�c�kQL�=��9�m���P�L]fV4ac�'\Ŀϰ-�F"w�=���V�ib���sڜ�Q�P�_W�$NS�:�Χ	�&�h�$`�?֪9�.��L��x�VxU��*Hz>����"�4mB��&���4U�"����W�0��*�w�9h�|��WdZ�e`��u}��?�-6��	y��!F�M^� �F�T섾������r�L�(䙪�?n2V�b�>��T,���}�t�]��_�J{_HE���,<Ua}ʑ�c�y�,d����D�*s��3}q�M.����"/<���??(+WK͚��_�	AV�� PG���~�Y�������p|E��$'�I�.S�C��;�/*0RZ���[�>�F�ϡ%K���-A�c4�4�H",1�� Ж�^�r��a�C�.ܓ�w�>�C3��6�BԠv�,��י��W���'��'�f2���Շ��PCF-�INIm$O_�KL�����'I��Y�Y����a������b�Y���Y�x�#s�s������Ӹ��/5�S����W߰�?��љ��[t:�L�ص����U�rdo.���ˍk+�|�;�i��܏<rȃ�m�e�2r�̗����-�d�p����������Ј����t�g�Vq4��# "L��P�vQR4�LT��=E$�(�A6��T�/+�U!������b�Dm����	Jh^�1��oNh��E�
8�Q��೴�:���쭝�ɯDGx(��cX:��g$?%Q%5X>|�`&���g�
Ў(|���Vj0M�O_�2Q�g�	�O�>L�UfZ������ɿr�#�ၯA����M�-3j�>q�OFk��˃�F��@���x�J�γy�Ҍ/�åz�i�|"ڧ��h���^������-�)�q0��}W�E�3�[�T7���Òzv�,/����*�F.9N��ʲ�Y0���Z!7���0�Ks=R� l͗����cn":2�QA:I(�,�y�i�^|�[7H��H'$�Y&�۪�b;��̅�R)r1�R��0X�3Q
ps��Pi� ���	.'��^�b��P�\O�h~I�ſ��f�3YL��T!*�`��_��2j��,ӛJ��|g�490�|�0w�ݮFX9��,��PN�)Ѡ�J�i�K������׉ZH�&F�Q�j�&��g�6u4�q��vr���SZ�Q�������y��e�J�\�y��n۽kg�_����`�Du�`:,h���6�i�ʹ��w ��i��pU���k�L���+��)�O=. �L���R��Oq��res}>��_;Ep#�pO�^·\�e׊�|��uR�5+�k�i�j� 6fhnr�.�=[�2LC��bn��Q0�[��L��>��CKDS� [�0a�$h2�Y}�x����nQ ��A9��I-S�#86P������0�`k:�`�+An�~�m���S�'����s�^E^-�*ӭqHs '0]3J�XJˉ����96i��x���6���K��>�Z��6�����H�3��E����p$���A�Ń
��K%��RU����-�S��
����,j&z�8� �q|����N�}\������A{�,��>Y��$���]�E��U�"�W��L,�/ob���nq�b�?�*t�4A�$���mc�$�`zE(�/�`��Dm�b��\((i4���<���ݓ��\��T�.�:� d`O/9Su��~k+J
������gw�ϼ6��8��5��8G�����$e��Y�$��M�M4�c�r�69V�V{��qi�p����幷n�W��t5��U0����T�ߡ}��Ar�3oK��cU�/#����i��2�jҥ�EB2�ad8?v~Hz�p�&��d���bp�eD
O���J-�o)����P�AfL���U��T��1��Щ�K{q
����"��2��^��)Xu�8
`�B"�`��(F��G�La}L����r�\:+�F���i3��l*s�q�1�H���:����#�Q��]<����I�Sh�u�ʤ<P�t�^GG��L�>�'oGnK?�?L��F�aQ1r5��i���j6����Y������,�O�?��˖�i"hR9C�1�����qa/���8xh���p��r1%6�=c��;ɕu1c���o��������y�t��=n�]A;�G�o�~�I�T�QY.$9��c�й	1�
}CL� .N��U3{#��lX�LfZ�]��W��K4F���9��KS
�6���F�1Z�'���'qDwqu* Dy�ȥ��ҎqH�QJ�^�<��R]G.w�W�O���Q����m&����� ;ڧ	���DX4ݙ\<n�Q��H����D�5
���]�2��Jk�Y�tE=�C;�X"�?1���1���LI+/~�N|"�s!���\�4�=���>�kp� ��E��ػ����:���tNw|�2"���qެ\R��nZx*ӳ��\���Q��{+�P��u^�x
`� ���b��)�:�6�	����Zp�M��`������ +�'�W��&�Ԓ��g��P09�s�ҽ<�)يt 3� *�!�cй ��]/�_�)Bs1%	��/��$0/1A,S�M�$_0��)Ss�1��@��o&h��5�D�;'��i�������Ot�F�%TT&�'����UbW��G�)Ϥ�0LSV��	��3F��dϾ�H"���&��.����lޫ��4�&X3z��샙���f[/��8���肧^�tܺ�N{��a��7����>��{Ls7'�1ʖ�(�b#���. l�ͫj���I<�.��\��M)
	���QYW9����b7�F�)��=�R�S���퀳���2�Xa&�ۢ`'hb��ۯ�o��B<��T'fC�F�L�����@HS�r�.ɭϧ�H�1�%+�& YT ��s�5�@��Nбer�έ��u��`�Ôx���앯|�@��X�q[Q�:�J/MQ�hI���(,�4ڠiBft�A.���]0[��˵Oy��>R{�ÿm�;��|��_?J=3�X�`	I������s��^��z�d�������cg��N,wiB.���Wc�20�+�#��;�'�6h��OfQ��O�����ĉ�O�j��nO�0s<Y��Оя��q�HL�-��,�Řaqc'��OJNL��Ms^���͈6��?��)�(9��<�͘��;�"���nZULz�Ҁ�ՙ�;��d��1R+�q�\0�l.��=
��&h����,w�q�#���ZK��ʌ��p-�vLX�J�^��b�$��|�\��������b�u��k�����5vR�''$��J�h��~�M���+�:��,(���%�����5Ls=3.}�S���ʂEurߛ�4�e�N���`[޵}��:tYa��� }7�76Q�}m�I-f�Ko1rp�pc����Rl�FI�w��"C�)��oc�&2v�L���uuz����*3X����<_:=�I�#'�߇�~�y��ͤ�t�������u.UPj��8�Py�ਭL*���:�B9�3"_$2}���E@@�����J����n���΍qŭ�g|��	�q�(m M_p����Kr��V%�'��Mg�T2W~G�I;)0�X0�����n��}��K�ݘ|�n�Qkt�jۘe�-����4����dɚ~#(�>pwa�r�v� �@�4$�G� ILW�w/��B�+�]5S��B {���7�Z�3o��-�짓�Qq���S	Ƕ�C��Ѩ�>�6�?���O}��?y��'��������7�~�C���@�U�഼!WX�������r�:벾s�^���/��w���T���]�ʿ��a	j�,���en��W9;��Egb:����]ź) �ks���͝��=�oXq�02��.��3x򦰥ʞ���������Ի�n�!l#Xt1��)����&!
��&2�6�>�/�τ��q�d�øC���T{�Y�F���)7��L�9?� @_B��*�J{\�<Hkb*
x0�A�������O�
rFбX��N�"n�t��o�&~����v��Bc�וK�-����N��z��3�l�'m��Sn����'F|�x��V�����OMl�<}���<��*�#4� ��/	�9�L�Ns�P�k7��s�Q�kZ�]��8��jz��LC��S�U3,&�+BKqY�`-�JsƔ��F���'��C��!�ޑR	����球w�Vr��`�*d�����0�@���e] ����E*!y�7!�*�2����'z�0���A��4�o�<��ai��\t��t&d]IP�Kֲ�6�n��JGȁ>�׼<�x�~��?������Dug8�n���߯����'6z�r�\������I̷T�	���g���,/]P��C�6�ϳ<j0��X\�O[�q�z}^)))�$�΄��K�O3�әv�vD	M@H�R�����>&��T5�(	�B_�Qk��Gm��HB�� 8y�钞�U�͎��TM�h%��KW`���ʒ���#����T�Ӂd�8���a��!_T��w�����-�\�&�L|jq�f��,(���R�3?ʂHM2�e�!��(��y��~��O)�;��*P:���;h�-�:W\֕�H�k��!�e�+1��yT(��@��.�֠SFFmE�OjCP��2�S�a�J��{Q��px�p���ns�0��ƅp���� 4C)+)��ehkGǀ'�B�H��x$�?�y`��� d�>��H#�0C�Y�3��bQ�W�N-͒�(�7�R�K]=�!�h5�G�ު�Jh�D:�FdmY@v�c]C;Cg�)�b,b�f���ʑ^�1�nd�����W�  �M�J� ˒�%Ҳ�,�V�I�v�Jh@�J.:�&'��r&����g3�<�s�Qr��"�����B�(:�cͮ/���Q��K�?��F����&I|�6r=�cr�edA�2�Ky�����)HВ�rb?�Q��很,Ƈs�|�Q̩O�)�@���jy.l�ɉ�[N���ɒ��6��������m�T��s�࿿��Ə}���+�o��|�ù:�۝R��n��-��<˱.�|�֖,�/ʪ�L���+�>uh�nsu�щUXM" �A&�}`=��N��0��a-t����n0|�.q`#M�R��%��Tۡ���t��4���� �#d��qm5���@\���5 ӺK<�p�`a�ƠD�JΏ�i7�K ZMC��*�aeҀ�����24\b�Odk�����^�s�wљ��!Y��NN�"�.�\�����1 `��h�]~|�J���9-�)�	���m��2�A�wQ��X�E+<�@ ���[���2�c�kl}RY蕽� � 42*����rj�b��L��zw
9&X�+*�������!�^,׽�BE�JA��)X'�������H�#,'�E�w�Z����9
m3���։�^�s����窢�\[�T�ǉ��^T���6a�T�Y!����'�/>�����@��C��V��UR5��0��� 
ڠԽ��'A�&h���RV������>Dd��К�0!Wo�Qf� ����.��� �'{Ke����fzz�G�IJ���k��
���e�cDJ+�r� �U
8�F��X j����e�}�@�����pT�D;wA�����#�S��O%��۪�ąu����O�~7΋��Ai8�UW9�AB��%�G P��9~~�/�x��[�_[�3��>��/��v���k��p��J�T�/��μU�eŎ�ｾ�H.���\z�ʾ&����MY��H���iB��?��vl���4e T�KQ�MZ�Z薖2h�=����6�HM#M z�N��(��p"���SB���IW�Z�T�Gֆ�x�PkW�-���O�+���h�G������j�$)g������e�BJó?\&m�"l��?ۅ3�X��r@����@6\_$%�x��� ʵc:��L{^��n�X��r54=�^�l�3��HOmf(�5�!��̯��J�]��b)-'Ȧ?C��;���x}50I����.�	��zAo�c�Xi }�{I�C CGp�?d�ڈ�s���4y�28���Ų���_�2��D��PpX=���H��u4{�qY::(��
9������E�L^j7L�#߁�/�'i&�+?
W���d�cH���|]�8}К@J�B1L4����ҭ��WA������Ai��
���hr1S��c���\��T}mA��ν�{a��ODjqx�^��[K��`=k#K=9�����%�z,*�/��1�=��3]O<`P�f��@��cH�@��]BO�iiczS�;f�
~i^V"�ecrxGHA���b�����!������X�<\,������MiH�D��P1�C�|�����;[�
U�I�#>�ʇ��E?����x�K;�q��o�|c�\#��d�Wѝ���9����_���Ӈ9V9���?�я���wOt&&?RLn��Vy�ߤ6Z�OyG�s�NKw�K��-���KK�*��I�k��}�h�S���B7�ͫr�QٰhX.��C��ʂ%0s�^�`Ǐ�よ10�'��J��}�rj�D^.Qm�S� �fk�]�ܙ�x�Z�Dd��0��a9{|H�n)���:[�gj�Ə���@�F���AqWy�l�Z��k��A�.C��M������S]�}��u]ڷpTJ�R\](KV+ ���O��M%��:�&���t�I�?&'�奾98A���T��t.�qY]�u�Y��H��������F��h7�&�&�:������>��
�9��� �]�:�vE���/���LH�
)
�� Kk��J`�e���R�g�^��0���N�t�?�kH:NG��+!�����4�_i�P�D-�9h�R~D88�X�����J1�5�d\]�/U5!���:��FDy�Pe���S �y�W���+���+��{����V��L�&5N��Z�@ߖZ�%ް,��Ȧ�^i^�H�!K��R�>xq S� �CQd��! |�t]�{<r����>�g����~~7_���!&P+`�|�o�G���y�鶚�M'h�=�	I��;�>/̳���q�򘬀fH��Y��}'����ܯ�
��� H���7^K����/޻����������S��O��⑟~�����O��'�(a�C�W�bI,�W�˴���e�6�Q,������������^��\{�
�'(��<+o��K�pQ�:��DS�i�H`�*�&�*#z�.?�%�=�
Ku)�B��D6�hu�^'�]��9չMV]S�N�vN�/�wD�l�#���8�T2kǠ���_f����EՌ�sIY]944eFIo��ep֬�Ȧ[H���I4!��q��V<>t���e��=S����4 +����Z:C5�� �M/�!��U;��� �<�������`�����Y��U�.�k)����l���&���6��Q).�IY5��*azvXb��{�����N0��j	Q/�rM�M����g��<*��I�:�2)Vp�s�Wm��1%� ��ͣ.���T&KW'd�������r&�*�HǺa�$VTl����'�#xt�? �7A�~)-���^�(e���:�O
%K�*ٮ��W�"*]�6U* �x�-����4�}9;��a��[�ў���ViL�-#R���\$ͫ���R�o�x��c�q�	��!�r���\^����]O�eC$$��M���q�m��%�0������o
$��~�O��*V0�{,Ao\9��#�IQI����`�Ͼ0���f	���P�L|��`��ftzZ���_�Y R₂����&�|�$����?8y���z�_�*8�w���_565�r��+���Q
���\8~z�~���MG��_��V���2�y�>fvy� �]"�rt��K̄�hU�m߃������@�)�κ/���Y���VR��t5�XԒx��ba�W��,U�����	@�ŰX��υ	��t�sϭ�T.�
w��
��{*��hR�)ޚ�џA��1��oe-|����D:��`i≝;�ѥ���Ta)Ys�"ɣ@� �ҳ�@���F�Hyb�3�<�!a�P�/��o.ɚ�4eR��*�u�<ʧiZ�C�TxgFt�d�b������=*O��a��F�W�0К�1��dHlţ��U�����F��&�h8��)e�Ʊ�W��e��b�6���y΃��)P��4�� �T�ҟ�Qy*�ʿQ�T8�v�*�R�Z��@P�`�u*�zD�q �j<Á6�$8<���WB@��!4/�J
��*��^�j4 �#e�I�eX? �c2�w�$��-C@����� ��)�3:n�Tc�<v��P/����܏��A�E��N-SR^(�4?�����	���A;"��5�燃v42��oN�ưf���2�VP^�H��j���>��Q��ׂ�b��O���X�>�AA8����H�G	�eY��<\��� n�l�/[�gE�=�-Z��}������P�V�	��C[b�kc^�3w�{9����>��e�,��#h�s7��+�c)��}�ۊ��sa����*���s%��jWڥ�Z�٠<}�!�Ita-Q�O��=R���Q�t�Ł[S���,p�L8����Z�8q&v�ч���p+�B�0��Q�>��s�r@ b�������5�A(��eGz���b�5J��&�D�lV_�|�x��ه�J��q��߽w��|*�L�����9� ZιޢBٶ� ɤ�M'��I��\����,ib3��(��H�ä'f�����7Z��5��s�2�pQ&*���)���a\�D~��n��t���!���a@D�N�8��B�4+P1
Jf��z:L6]���e��q�U�2/L5MNh]�H���Ba4�Ӳ��H8��ގ��B���S���W���ӣ����e���:�IP�)�d�j��P��Wsx%A'xp
��+���o��<�`WQLw:r��w	^i~���	~Ax=�)3V!�������Om��׸��/�?�2i��0������TQ��@ets�}���$F�>�6e?}������NȺ'�g��� 	��S����f�ޒ)�)��Jo
���s� r!ꣿ�L��v�aLn�w5gM������9��ƥ��5f5��cT�R�(r�t@α�\ra����oG$���~`�H'U� ��
�TΉ��q�2򔤸gQ��i5w��,�2jη� �1�>�e���jQ��*�Z&�`IͻBh�G�a�B;�� ����j	�#r���RW׏H�Ż��S�	�-"pr��X�=
��,���cM	��)�\�L?�F�JSA�HwGX����G�,�A|qY�Wڼԇ��ػ�<�Y�S�&|�l�6��Q6���`�*JD���"x�4��vA���RP1���W�fIx*$�D�i*ǜ�3��4X.�h*��7߾0'Go����Lz�ʸ7��e�o�٧��ĥ�yB#0����.�tt�6���a��ऋM=��$Ï
Z��U�Ul�M���Zi?��ƻȗ�O�2����p�S��t䁟T,�ր)Y �n��bÆ�o�'�2��'>�p �����I��dT!��/8�^�����%P%G��p@(擒�k3����.�Ed��be�7)}	>$~[ PW��^��zD"C�m��oL�@�䋶�7�e�∄0O�� L	����I�+Gh4"�l�8�����8�C�d��t�]v�l�eJh�1�R�Y-��Jp��v��*�Á|k���g�UB���J;�5�'G�f0���ԔQ*�\3%+��m��/��J�B�Tԥ�S��u4 �Q��`�3|1��zD|�hqWЍkN���գ�2u��M�����a9
?�aCSj]t*���36}=�TQ3�c� 4eYX�\W!��*����^��,���:�_��nsU�6`n�g��D�#��%�.��ۢ.�@� �n7�L���"�����%�Q�I����S<e���+�qY^�ū�R	`ˀ�i�x��
��|���4XI-G���������e���������N�<��1��܊�(���$	��^Y�� B��fz�R{�s�r.��d���r�<��ß�����wy���m��3�LfH���p�2h&w��6��:ᔽ@�օLq�ºp���Џ6i�����a pKȱq��aD��u��i�&?�%J#L���r�WM��Z���ȋ��Ew�_r���el�$�m26r^q�Eif�&�I�6K� �1h+_�z) `��N�g�g�x������E��n�n0M����I� �r~N۳�N����`�mU ���d܊{���@ �Rj�W@��b�
� ��NAПS<�a�AW�D\Y�S�{`��ß�'p2�6D�K�-O,<�S=K.�%��ZP��ك��t���h�-hj��@#��i��vD��B8�#��7D�վ8KזK�"��||X�D��A��Tld3'�:�L������|�.A����ٚ�υZ'Cq��p:���;e,��$����}׼��Z �χ�,�QBЊ��mŹP�K��X�C6�i������E����V�e��㍥�.����8�9��8���hY��#��BH��Ls$E��	�	�e
v2���}���F�v�`���i�K�o�~K���*�&�0��(��7�N�w.]q/|D�1��˨�͝�[�ܲ�B&�y!�Q兟:8�:��U�NQ@��X Mh�� -��~Y��U5�Kh�-���P�e
�f,x^!4|�`�A��{^6^ݤ򫱭|Ω#1qC����1?I����t��U�ԻC��n� ��cȨ� �RGQ�U*1�Y8n��ݾ�Z��&�8pȡ�Ay����G?��R�����3V�� ��+�\��W�B&5.xc���py�SZV�%70�i $�^O�٤6�`�ccC����G��{�l�"ٺu���|NQ�t�G�Fdpt�G�)�>F���d`I�	@�z�T/(��W�
��u�pX��T9�!ҵ�fh�.��=����?�0=�)������<U����k����Z��V��s������0@[BB�`&u��= +Qƈ��/^���|'��������h��d�u��H�{a����~��@�{ɴZ����3�H¿��4B�4:`�Kd?{�]���� \�4�]w�m�s:W��`���&�|��cd�uP�H!�"Ӷ� S�3��M�_ Ν%ހ�4C�����y��W�v��l���$������Z��W@�D{�9D�,B5���H�_�F�B�D�$��h��<4����6����h�G���)>U u+'K֚�:��(� �5��4"�� ��v��w�+��l��A�TV�t�]������`i��i�]�vB���Yn� �n�E���0����ft5�����2����+7�騵��R-�_s|VCC�����B Gu ���,e+�� q�¤�=���ڤs�
&J:)O�4*f�0i2�-M�9��;�h���1�0s����q�s�Zh��!`K�5Q�����W������(��gf>���%+�>����k�����}���C��VQ�h2���-�l"ý�TL�c	�W��%>��������ۉ����lk�R���r'�������OqZ�FЯq�%F�$�f�KS�3 ���3�:�?��3�!�P5����~Brs9,;�Fh��D:��0��� �Vm&��kȣ�>�2��( a�0[��!�ow����
'��Rk�䁲�i,��� >4��P���IFK��r��A�T����G)NM7<���e��<��n灤��z�]��|�j4��4�<`�F�]���4幺h�/��`KوT��y16aS�R�T��_�(�v�¦X�Cw����"�%K��3
O[u0M�,t*��kQY��#<q0.���/|{-']������ٳ]���������"����$q�J:�LB���H�� ��AC��$0�v�lRMH3�����yRn�N�b+���s+v�%hM�
7�$��a���EUαܪK�ʆ�j���Z�P��Pռǵ����k- }��=2̛�Aa��vP>�A2	�"|�&<��)���nR�)U���<�+if�Se��/j9@He�����f��9Ӊ�i
�^୺��A�=1�[�#菥#�L"�Bٺ�P�[��s䙅 ��HSv�}WN��δ��O�M&~��j�y�2y�/	�YʞT� 넀��l1hW�:�dA��|��T&�}�2k>�;yh�#�m��	��d#*�8�O����q`rN�g>�Z�@(`���c  �5��d��d9q�L2X���vh��Kg��5�K�g�us�=�xx�,�}���א��g��W���(}�
:�~!�n��S�*��b�� �&�R�5�ͱU䣊��)� � �;�_ץ**�3>�{�5M�}���fҎ�wי<e��K�3��L �җ�LI1���Kj'�8�:�EJ������Q�r��y����ɩo
�1:Z.����\��4P�R-sj�R�U��PP�!l��v�$�S?��&���3y��nA4�Po�5�Z ����Gf�%l�Wn����Q�Cc�̆��n��Woo7�];NR�DR�~���æ�؋�)��rk[�>W�����yA{�䚺�u������M��}Z�
�:8@�
!]�xVh�R9_4�Py�	Q�I��f%� <������AK�c~ep��d��M����	�9:����^�Q/�B֒jO���8i�丣����G�܌kC��<m���)}}}���/�]���k�:偧�QUR��ٷԆi���7�	WV�7��9:�c�1`^ʲ��f��N�><{�Z;�qq��,lo~���*\;L���j�Nկ�`P��:��ʔ����p�Oy���C�C5����`ᔜ*v�>k4;��qjY�Ǳ��s��[:!q%0�'56�3�.�k4�R�e5��7�zy���L3�����io)\�յ^�jK�\g)|������,�YjU�N�\��44�T6imm�9���CГ�#{aVqÝNj&�_r��!���-���,4��/l'���1ddrC�@dL��ٽg?���{���FG�i�B�T��%4��c�Tr�l��>�/9�X(�:���/��~�N��$J�V D�jQ�W 	']���U�����Y�þ@[�W~���d{Ք�s��8)��ߏ��s
N���K�Hg1�T���y�b4!�tV�y�����n�ﺍ.��U`�Fڋq�JR=��W4c��k4�5z`�O�z�ٽ�4�8���T3�M7\g�W���!� O�E!_���&�������}j����ݳSε�V�Ik��12~���5ʡ%�lU�'-M�M���f�
��~o�
:�[@<\��ܴ�<�=�دd���u'O��D� ��D9t�ze�.�an�ٵk������ϡzzF�ԉ�$x�|���{�Bp��~J���"�B����.��k\S6����<`�WtQ�ZO���T|^������Wm]���>t�g���l���_Ǵ�L��0i嫐a?1�ꙺb|c�������%mm�������PN=h�)-�On��Mq���i%�k���`.y�T�/��a�
�Nѧδ˾��d���9�Ѽ�宀i����':$3gs�)_
��4X7�C�z���? ���t�+9r�P��E�����Ν{Qϸ���x�i%S�xΕg��P{�I���,e�r����C���_�� 
iI�ʡ��N�18�4��Zi��� r��m2��n�δ ��==��~���Gʥp�ɏe��;��懚�ԅ2s�Q�&:���HH��1jj�0}4�9�>�i{{�|��_@�����o�T�e�0��!����|���$��M�����O�8��M�	�=����.�  .fIDAT�cy�#0�S���%a�������u�A�S���B�l���L2��1�a��+����M%~Q�M*���U�l}iF�Y���|S6�^�S�|i�侀h϶[�.��i|�=�"��{��g[����>=�EL�Ӭ�ӟpk�Qujc�i�M���|�[ߔ/}�8�2;��n�W;��1����͏����dc��D�'��A��?!#}Ǥ��f��G�`:v����'O�&P��H	N��
-�,�wSS-���Ǩ���2�V������a���(۸s����?-��0�P��y��3X�s�\���x�'���!h9�My��������R_W�x�Rp1�.�A�d�Ag������~��[x�<�I��;e��η�?��_�'>��h��2�{�c8�G����|�A޴�j�*3�R���#s ��N!h"p?wia��hI����?����砱��(s����?��<������P�ot�����WgA&��l)r��� Y-ӭ<���S�_�`��G�쓞�^eB��'&I�0��~������~�l�R�t�^���)p��=z���ռ3���*pn]��ǏSگ���wˮ����c��Ҵ�&i�'H�B�ZO'��dD�Z]�!_�~��^Y��,��5��������e6����s���	��v��Ӓ�������������W`]<mS�D�7��'�|^Zc
x�<@ �߿_���/�A��Ka�mj��p�����Pm�z�Rڞ	��2�Ͷt�ڸ�|�	��W�2�Pb�4��d���HwW�Ť�6#f�C7�����<d OɥH����D�%�*���w���/��7��ǧ����� tY+��ΝƦY��Q~��w�3u;�O?�����_�����ʲ%�Ngv%�(5mٺ-�\0 vx����3�'���KO�;,�V͕�K�V�W��E�я<鼧ޞ=�����!L����3�B�T��J���y��bC�E9�̙����"����gD��L�E� ?�w���B��d��_��|���Y�t|�/[�$���Ǟ Xʕ��N�&eE^³��8��� y�|�S�T�I�}D�5��?�o����ϥ�l+ �6�2�c����aH����{ArQ���&���a�����Jꚕ����]�h~��d����^z	|K!����Ȯ�;�Y��F�'R�4�-����1M�qh���6ǣ�j`�$�e�����ev�
�K�mX^�g���U/�v��2�����.Fd�#���{AowH��7`��n8W�� ��̴>�dW��JK@�X�D�HI����N��׿*�JCÂ�U�Ba���AhyH�C+e�W�8����f�c��͎D�qPd$�5����y�1���<��;d�ҥ�ɍ򩧞�_��q��嵯}M��9.����1�ڭ<f�ڗ���,[��f�&1�/�������F֯_/�W�Y�B����Y�s��硵!�ͷ�KI��q�3��Ӓ|j�PC��҄�e�k+dq�Ryq��|�[ߒ��z��� �ʓ���@~��O~��� g�*��������Ktٲ+>y��ڿ��fϏ!�?�Bfa�������w|]>���D�<����i!����m<���<��I7���)e�.��ښr��D���Ă� ������nK`�?Y  )���t�+�7���|�3�E��)���륮�d�Ai�h�0�O<��$`v���S1̐��	�AKZ
5�J���&)m��NG�d�Ѱԁ����ԦVU����3��W�E$�R5Ǩ���ꖗ_~I�Z;��w�%�kICJ#��'�#� m(�g�>x�'�+�GhQ��q�����U��>"O=��4/n���
�#P�9r�I6r2[k5�>���v����)ߘd�����G�J�vE��y:]�dr��������+���-k*��|�����7�Lsѫ�_����d빾����z& ]�N��D���S�&	���t�F�4�@)��a�
��Ϋ�k_�������W�&{�����˚5뵐�-��ڋ�����.&�����&\�T�l_y��C�����LFa���@&�!&]��Rhn���y�����dh8$���y��q������ $˗)R�~��~�'���@�E|���F[�Pj�CS�P?�KD�D$s���Y���!��6�2�6���H�7.��ׯ�#G���f����3�OV�^zN��ʴԁP�~���\�~����;��jR����Ȝ18��a�0ߍ[��"������2��O�ܰ>Cya�Kr��� �/�0��WV ��B�N�MgG���;����y�[o���48������G���m������`P�L��=���>�c��� ���+��������c�O?,���/|�s�E`�F"t���R�]16p>���5�b�" 9�vF��ag��}`�W�%Y�:�i�aӇ����%�8�5����[�"��' ���HeY)�AHsa5��Y(�������wȺu-�@�a|/R��߫i?�ɠ���������F���}�_�0�^�����/�T~��_���o�/G�f\����DA������;��;�V>uf!�>����J}������g����Wj��d�����(?1�OyE��ş�+���G��G��ة�4�C�6*���/�C~L�w��L���X �����L��VCe�C��ұ\��V�8�����j������ǁu0��j̙Y
���b_A�-�����ݷ����i!V������WL�橓�nJ��x�!�C~����#�A�Bf�熄$�P[���
�����3�S/6I�o��=���ߋ��LP�c�Ǳ������_/���[�wQ��������,�;N����;Z�HiN��ѧ�j�4^HrxwHqFQ+ �M׮����.�ܧ�­m�0/�k����E�cL0�A�# f��z��}��r�=[�kZ�UV�A93P(C�4P)F�(�,��p�a
�a05B ��ʫ�m��@ʁw�П=����=��A���>'/�c��C7ޭ��#�{���ݿ�:�5t���Ƚ6��GG�$��@/oM*:+��c�o�ʫק���W@Um]#��"�������d@
N���e���0]���07�����{�*� O F�RG��9�KWf^��|
�x�bv9�P(,��	+�@}��w�h��~�7Jj���ÇZ.���d����ЛnS�1�O\�yf*���a��9LRˋ�j
��Q��9��)UЌ��@b��jy���&f������m�1�Wk���!BC	,|��|�[o�?���!!I���8����Ag�t��&�?g��|K=�H_��\�sT��Hѷ��������.�kS���>�{F�>4�s�ur����o�K�m��E�ԁ��C��[�;G�'R�3�z|�	�Ol �g��1�5����5-����[h�v���4Ҵ�T{��/�\aCT�Co�Uފ�a�����>qY�?�ގ!9<R��E�^��;D�AoL< [�d>K��y�`2��g�쩃8T��<�zm�k��̇� ާ1�yw����LpѦڒ��y��߿{s��>���e�r�n��n�<A����i�l�sǢ�W�ڌ�r�Z�����������^��a�]���҇��w_#��c��T��9��kF�(`�|0��l�*��$Z m$s�����B~+M��1�3�#�N<�/������G�7�TCȻ�L�ԷlY!��f�Md&��4�O{�c�99l`�i>\�˕k�R�!�?�����~�<��`*I+��lY�|�����sς
����7ܕͭ�	�̢%u�������8I�04����}І0�An�s����Ά���Z��Q9�#"Wos�||
H�����;aު��������DmT0 ��C�.YZ/���塇nQB�Ԃot��TQ�T�ҝ'Xb�	{�<�`��xLz;�r��}�+Ђ��1����*�8�K���5��D��,\XX���M���C�19{,"�C>i|r�B�.)�	O@����kN�͘����B����,?��G�3��#ٱ��#*2S��I��0����o[����**�4l��	#|���_T��<������},� 7ot#���d�n^� ���B�I~��S��u�=����\�k+�ȍ�g?F���$�|z��\@��S�jq�y����ˢx��8��N�du�(k�.�(���k��Fhn����#�d�K�a*(�acc�����]$��DH����t*��N��İGz�;f�(��Dro�3H2�3�\�e�643G�e�;�Ӈc*8���'�Z̗0ۗ�F6�	z���H�\\�����Fn�'��wsߐܥ�ܷe�	s���)��@D�Ͼ���$C3��R��e���(��c�>��-`En��|��r�h�ڬ��R�ıQ6�_>����s����X��Q��i�ʹ����G�>��7��И�<�kn��]�ē�y�>�����@~��3��R��,´�0�韾���+��+���`_\���̅9/QN���0�S���d>wKe�s��XF������?,o~��ʳO��A��W����G?�y��7+�IF�j($����Q�r��N�]���h�n����!ܕo�aU�>Hr�M�c��~y�W��g�zL��;�ZZ_Y�q����ɖ�+aV���~��{Q�;�
������2AD�b0p'�H����Ϝgn����OG�\�^��͝��Z�/t��X����!7n�
s3����l߅�.]H�� ��A�Ms5�!�Jl�˵6p3���t�0Ik�I��+�Ç��?�#��:[��N��ƭ ���5�������O�}����F|�{ $���Cr��\�{D��G^?�Uk�\�|���J���m��[�W�2��+�� �_�݊(�N�\��S���X���ئ	��<����u�_8�)�����	q�⧲�\���[�-�)i��o����_i���19��A2�0��Z� �i�j���|��EМ�� �U������̀���J[��𩢶�J-ԘB���576��5[ƽ������w�eP�4�虷��q��Kn�	c��v}�	O;K����$��.���v��R����g���k�C�p�:�k� �&�H��	�ڊ1�?�D�i$�T,lp�Ny9P�g!4"2�뒒����8�(���o�w�����l��#HwQ"U�P_s����f����v"�p� �E@�&L��o���Cu΅ ��$�(X���rd�S��f$�{�x��:��A�~��}����V����O��؂�F,Y���S1�_Cm`�Z��>�|�Lk:#�Οtʂ%6� n���5�ٿ\x�F�5i�`X�C�g65V,���Ѕ)���>��;��a�˰OIK0's��#�+.���ɔ��P�a�\��A���;�a"�d\����U*-�5R���vtC�t~K�����IK�a��7�[τ�I �F�����"��o(�7��:5_\�Kjvb b�
f���?!�p� �Q��p��A!O�k!��"�5�q�,�ƔS�-&rMG���~Rg��၄�j�Q1@tp���L��Q�����%��j'|���ԈPzZ��c�`T������P̰g�.pԏ�W>K�%2YBA�2��8;�Ťf��`�����z8�4%�=ǡ�=qR�^x؋�h��N[�8�n�V|w� ��b��oY�/&Xb��Ӵ��T\�F���g耀������b��5������%���r+"LtbI3Y;f��Gg��;�����)."'z�d� ��P��#�XM*$hT"�6�3\ w��*樴���q��:k�m7�W��2����v��O����;~J�=r�;(Ot� �"�l�U�sDxV�^E:^�B~���=�&z���ip�~b�ԪU�U�]�u����5��J�ȍ~&��{"r��/Ƭ3n��+�Z.�/�q�f$��R�3H���Je�|���Tee^YTX��jc���:��]�@��ː�i��p�r����F�)4{C҄����~�"�#�U[���أ(4�ѣǠ���d���u�y��@�D �q��S=��Q�����>�<�Ѷ�ᑦ�p����Z���hfĖ��ė<�[�#-�Vڌ���I �Rj�fRx;����x�k�+�&��:'�v�7K6�-u�K{��y��3�Ox2��|��C#n)n+7��h��r�[�-�p��p�s����܏R" \^�ʱ�腦v�P)̓��s{�KX �0�������=��^Yc�aIxW�-,�V��p�������� �x���7��1�"�KϘ9�g2��^N_�� ���l���'����y�c�|�<`��}~)�xIt��L�؀���ɶ���=��%px�#(E�\� ����/�@�q�1���"�}x�.'BEy�%s ����b�|ȍ���@�!S}	X͓��'c��+3F�d�:�߈
�lP������zIxBb�_}���l�^H��� M����q�LȢ�.�_�U�\�c3U��9�=-�!��v�eW�
���Jw� ޟ��N8�G��O�l����'h�/xjր#���㎍Ri�Z��>y:,;��pևVq�����쏻���X!|T���;�
 @J�4Q`j�[��+m������93q_GL���t�G13!j��6��|�kdy�H��JF[\S����}�����v{VD�������)8Nx���8اm2�8��vw�+K������v����Q�F���~mM<|k}�cr��0�������Hg�H����}� �u�[j�)-���0]�d#���TEOJ[���74�z~���_��#8xKϨ&����9C���!Ҥ�L�y�s}�4;Z��M��cv�Ǜ���D�@�ɾd��d���!�y�K���+.����LF�r?+�8ݽe���-�x��M��7���y�t:�?��� &�7�YB8>?R.6DC�=B:�,�i�9�T�]��O9w�$�&��4���N�݈�3%�:����"���w9��G~���
\҅�w�J����[�S�!c<������Ծ�
V�܁��7�I[_�v��O.e�>I�&D"Ec.	�ȉÈ��#�-.E7@Q�) Oi!(L!�/�l����:���l�����g����YRR���n�6AÖ�qʒ�vP�)s��@������c-"��sr*P
�.�Y K�Of�aB�$�֧�R��~�FZ�k�y5F]�ı#�g�� ��iBٷ���(���?��K������Y�>c�2�J'8�����f�n�3�wՈ�asٷ�G
ޮ�Xo��G��F��+R��8�OEf9���>��! �cA�p�h	�4M�3�S�oZfS�(� �"�:& ��2������6�����쀥�9�>E;Nì&����  ��q���\W�ͨ��x�8fk��;a�<�J[T*ԎO2���g'\	�r=�mb����=�������9�Ꝫ���EP�l����܋��-�8�V..��7ܼ���]]5|�۝��}�[9���� �˔���$_��|č�'����н��'�Jrʫ��p�j����oiM�6s�?��h�b:q �h����rhB@6�OC&��0�)�?U�;O�I��[�#�{����C7� �Hw$0�٢��B�A7 �ߕ�rΕ�]�7S�l4����)�fGX��zT�n�t$&�W��(5:41�����SnR���ME�8����Jz'	I�{'a����.���Σ�3a&f]�3��ǂb��'���������W��C�b��ahpZA��*��h�'�h�b���vP]�dl�HA���0*/�:�̯	̟���_��
�Y�,Ml��-�.i�ig+���|�1y�:����$a��@����?
(�&�Gq�p��: F|hgh��2�oo���I_!r����ՙCH3�}@[���
RG�џ���iK�bnr���짶c�aͶ�������SA�?����4\hOZ���P`&�	ڊz��۩�8hҨ��9�%�6���5�C� ����,�ר���7z����}�5_��ln�3�k0͠�['Y�X�@<1drN�4��ųi���w�s#����/�v�b��/ˮr+SsdQ�ZV��@���
���y� ��i�`�^N�F0GP4�E�'��'�K�Жb���1 �����E��ʱ�Z�_4	{_�����2D�@���."'4K<��Aћ<T��F�D-p��ȁA9�E-ni����an�|~hl�<�6!����UjG� 2��e����x_�� W!2�l�_¯�y���F$�	��(h&�P9��Oa���lw-#B�,�`��V��Q8n?�_A��lk�;�'���9����>�ep�p��͕��z`� �*��|���
���OF ��Q���������V��cpX?߲h'���"8� L�O�I�ݲ"8ʣ��hb`D_�}B	�ta.ӄEߞ��(��4�#��>��R9�"1J�h��x��ȧ3K*;F�]@4i/�
ƪEb���yD�}��b�OS�wg��@����YzTm�.�gn>������5+�?^[�;򶻛{/N+r{�\���Z1�\��$�K��*i~ip K���*PQ}Q2+]&�Y��`��P��""�iN�����,u����Q�B2��<&�QT��(#���"�6�	"� [4�6���D�al��d�B�S��~,�ϷK�	���ŕz��b'�s9+�c����
�Jo ?%B��(L~ a��9�0g���upCN��G�� �5�_(=�A9���c���`���n��޸G��.��пf6|l���b;G_p���J98�����Q��D�s \B�돂�%j�T8�L��h�]?�	0�����c�`�*@���;Ɋ�~����>k��Bĭ��</B3�V��pn�7�1m��9�EQ��(�w  }���>{���
����9v�L.�ÆA�0�h���jq����)�É�N�Yw�Ă2�$9�6�q5F�
�H�s	h�Ƌ�Wj!2�\��C���s���r��a�p�#k�K�܋��qC�H�9�
g�v���MB@�(�w�*+��ݴ�����ߛ�g�Vu�i�z��'���'��r%staS5�׬�u�(��9j� x�Z��@P�F�ĨRxۤN�5���;
�h��6�� $ �
m !�\`�<�o�\��D!�� ��(U.5��gWa�<�����T?@��x�&M/�@H��Ɛ�w�c��B5�U���"��Z��GQ��3z��Z�Qi�Yȁ�`���C��T�!@�*zY�3�ᛕ�f��qګ����@��#`������Ȭ�� �4�؅�Ƒ&���x:�q��F��J��v�����M��uE��Mn�J&l������ �N�җ�'�[o�?�J�+�ť7V����5~��=�W%�v�"�2i�#QJ_>$�.±�Jh
��V��o��X��c?M�*6�K1/'{u�����ٱ�����-_X�����/W�d��<`�ػ���2�?���iA��X�\��~��`輵(7X��D�O���o
eZ�kZ=BAj��M�rP��2��X�v��E�8!�/�QA.����,�%�?f�#ᚪ^8Z��1���}UP�SId2k1�[�թ����#�H����9�4�z�P�.h�aی*��T����P�Og�fk
����n�� �ߜLʟLM�K���75}�&r�����h'[A�6�������xy�R��n���֤��1A����#Od��P��Q�zච�_�&�$����qfþ0�0�(uO�B��Υ�=����&V�G����E^��k����{_��H�u\����a�K��/*i'~]�dH#�3�I���HT�I吨�&&b��tO���U�HuPOތ_Ȓ�j��Z�?F�!ʥL��1M��.'EJSB�R.
ͥ�S]��ժ����gZ��oj���*�{���E�@rR�u�� 3�mL|���ß�V.E�i��u>
�?P�0��|'`B��[�3/N1������>8�#�� LT*r�����\]�}b����qOK�W/N�f�)�iV�󲬌�7-�ICe�����nX:O�ih��~!
��S�P�(����(U�L,n+i�L�>E�=˫\� �v���fg�w7�5�vk&�7�|������#��ϝ��L�� ʔP��QUJA)��$�����a�$Y�f����s�LBp��T?�ʀWJwLw�LN��A��N�|������pf���&$�va��L�r���/7V�,]X��r���e�r���<`���0�7H����<f���{���QD��cN0�E�^��]���~�1�ƪ]�-������� B3mӥ�?7蘡uӾq�o:���'�.�2�M�~e����x^J�����~��n���V����P,�ߙ7�G�<d*��G"3S�YWz���}I�1�+K��ۤ7���[�����Z���p ^���֬��<H���X�ʫ�Q��f��]9<�"ζp�_P��R�����3N;2�i��22%<��e �w'X8��[���e�<��qwt* o��ZA�?�*��=�Ku�p�����s��;���A����ebY��J�=�%��<����W���:���eY4��)�/���u/M�ʨ������o��t*�K;lϩ�7����[&�W���po�J��G������~R��í�R?�?T:ҝ��������Uah
eG(A`%���z���B��8 �FKR����T�  	�'�q�d�J`�/TfUT��a�Y�OyG�Z~�� �b>�����0h�'����me��{Y�(N�a�Æ0�d?[�l
:68Y�rs����!�N�P4�����l�|٨�i�_s|������~��8�{��=�ٯ�q5�꒿���a�)B��.dTa��bo�/9�C��������>�]3�R�:�3=2-��U��'"�p/Ĳ�l��NS��0��[�b��Н�_]��L���/γy� ��2,�틠;��D:���-$e˷�h�|��>e�̣%a��째W�H��+]p�l���N�R6z�]�Ek�O��"�=bل�u�,�q���h?J��rّWQ�����b|M��q�o^�	s��i�� $�'N̤������u;���n�kN>��SuRE?����"�sٺ�v����)]�)!h���(D^�}a�/V�b��	> ��;������*�<�����=0��=`�y��ʟ���}�
q�lk28D�� ���BJ5�e:6Y��G>��1����z	ճ�d/	Y�:�3ZB	c-��8��9l�C�� M�"�,��$�����G�N��Y�O���U\�*s
o�y6w��Tߛ $�-`Y�q��3ԩ�)���|7*�����U�Ӕ�C^W!\3S�Y�8@�� �į�����S���[O��Ɖ����;�/Ma���6��=0�����Z������    IEND�B`�PK   *�4Wt�؈�  �     jsons/user_defined.json��_o�0ſ
⩓����e���5�T�n�M��ƟUU��>��i7C��{�����ٮ�
aO��Dld&{b�e%�L= .p�Z��u[Z����/?.�������*�h-e&Ui��>/�T�}��V𗻚�2Q�2�a�9x�3'�>pg���3��N��)Qť,�����}��@�[d�����"�����Κ�@VE=��Tmӆ��}L�*{}v�?c���=b(M&5j�l��u)_�^[�W��t)S����~&�PW!@[#�Y��K����4Z�]�����I7j|�>��Hz�H�s�g�����Ы�i*��
R*��_k*�\[g��s��D���ߋ�5<7��@/�jx����M� ;b������a/���@��ˠ�m���)_�Ӌ��A�Ҿ�F�?uGSSz�`vd����i}vqDCw37ո�֏�}��	�7������>ce��l��ʼe-wiچb�g���N�o
/��
E)��Zd�(7Q,�Y껵̓&C�cC�O�i'��^'�70�x��'d���lF�Eqԕ��� �/�a4#�r�(�@ໄa��G�I,��������x��,����;�w<xG������z�BHG���x���ވxݧ��ם
Ɉxݫ������xr*]7��Q�d�n��|.�_pr��]p0���fp�oW�?PK
   *�4Wku��"  Gb                  cirkitFile.jsonPK
   Є4WUo�H̒ �� /             �"  images/448c166d-0905-4b6c-8bbe-acf1d9153e5c.pngPK
   $�4W�'TO/ �. /             е images/7789289e-5858-4b68-a160-e98940e09304.pngPK
   *�4Wt�؈�  �               6� jsons/user_defined.jsonPK      <  %�   